// --------------------------------------------------------------------
// IP_HELLO_WORLD_ROM
// --------------------------------------------------------------------

module ip_hello_world_rom (
	input			clk,
	input			n_cs,
	input			n_rd,
	input	[13:0]	address,
	output	[7:0]	rdata,
	output			rdata_en
);
	reg		[7:0]	ff_rdata;
	reg				ff_rdata_en;

	always @( posedge clk ) begin
		if( !n_cs && !n_rd ) begin
			case( address )
			14'd0: ff_rdata <= 8'hF3;
			14'd1: ff_rdata <= 8'hC3;
			14'd2: ff_rdata <= 8'h00;
			14'd3: ff_rdata <= 8'h01;
			14'd4: ff_rdata <= 8'h00;
			14'd5: ff_rdata <= 8'h00;
			14'd6: ff_rdata <= 8'h00;
			14'd7: ff_rdata <= 8'h00;
			14'd8: ff_rdata <= 8'h00;
			14'd9: ff_rdata <= 8'h00;
			14'd10: ff_rdata <= 8'h00;
			14'd11: ff_rdata <= 8'h00;
			14'd12: ff_rdata <= 8'h00;
			14'd13: ff_rdata <= 8'h00;
			14'd14: ff_rdata <= 8'h00;
			14'd15: ff_rdata <= 8'h00;
			14'd16: ff_rdata <= 8'h00;
			14'd17: ff_rdata <= 8'h00;
			14'd18: ff_rdata <= 8'h00;
			14'd19: ff_rdata <= 8'h00;
			14'd20: ff_rdata <= 8'h00;
			14'd21: ff_rdata <= 8'h00;
			14'd22: ff_rdata <= 8'h00;
			14'd23: ff_rdata <= 8'h00;
			14'd24: ff_rdata <= 8'h00;
			14'd25: ff_rdata <= 8'h00;
			14'd26: ff_rdata <= 8'h00;
			14'd27: ff_rdata <= 8'h00;
			14'd28: ff_rdata <= 8'h00;
			14'd29: ff_rdata <= 8'h00;
			14'd30: ff_rdata <= 8'h00;
			14'd31: ff_rdata <= 8'h00;
			14'd32: ff_rdata <= 8'h00;
			14'd33: ff_rdata <= 8'h00;
			14'd34: ff_rdata <= 8'h00;
			14'd35: ff_rdata <= 8'h00;
			14'd36: ff_rdata <= 8'h00;
			14'd37: ff_rdata <= 8'h00;
			14'd38: ff_rdata <= 8'h00;
			14'd39: ff_rdata <= 8'h00;
			14'd40: ff_rdata <= 8'h00;
			14'd41: ff_rdata <= 8'h00;
			14'd42: ff_rdata <= 8'h00;
			14'd43: ff_rdata <= 8'h00;
			14'd44: ff_rdata <= 8'h00;
			14'd45: ff_rdata <= 8'h00;
			14'd46: ff_rdata <= 8'h00;
			14'd47: ff_rdata <= 8'h00;
			14'd48: ff_rdata <= 8'h00;
			14'd49: ff_rdata <= 8'h00;
			14'd50: ff_rdata <= 8'h00;
			14'd51: ff_rdata <= 8'h00;
			14'd52: ff_rdata <= 8'h00;
			14'd53: ff_rdata <= 8'h00;
			14'd54: ff_rdata <= 8'h00;
			14'd55: ff_rdata <= 8'h00;
			14'd56: ff_rdata <= 8'h00;
			14'd57: ff_rdata <= 8'h00;
			14'd58: ff_rdata <= 8'h00;
			14'd59: ff_rdata <= 8'h00;
			14'd60: ff_rdata <= 8'h00;
			14'd61: ff_rdata <= 8'h00;
			14'd62: ff_rdata <= 8'h00;
			14'd63: ff_rdata <= 8'h00;
			14'd64: ff_rdata <= 8'h00;
			14'd65: ff_rdata <= 8'h00;
			14'd66: ff_rdata <= 8'h00;
			14'd67: ff_rdata <= 8'h00;
			14'd68: ff_rdata <= 8'h00;
			14'd69: ff_rdata <= 8'h00;
			14'd70: ff_rdata <= 8'h00;
			14'd71: ff_rdata <= 8'h00;
			14'd72: ff_rdata <= 8'h00;
			14'd73: ff_rdata <= 8'h00;
			14'd74: ff_rdata <= 8'h00;
			14'd75: ff_rdata <= 8'h00;
			14'd76: ff_rdata <= 8'h00;
			14'd77: ff_rdata <= 8'h00;
			14'd78: ff_rdata <= 8'h00;
			14'd79: ff_rdata <= 8'h00;
			14'd80: ff_rdata <= 8'h00;
			14'd81: ff_rdata <= 8'h00;
			14'd82: ff_rdata <= 8'h00;
			14'd83: ff_rdata <= 8'h00;
			14'd84: ff_rdata <= 8'h00;
			14'd85: ff_rdata <= 8'h00;
			14'd86: ff_rdata <= 8'h00;
			14'd87: ff_rdata <= 8'h00;
			14'd88: ff_rdata <= 8'h00;
			14'd89: ff_rdata <= 8'h00;
			14'd90: ff_rdata <= 8'h00;
			14'd91: ff_rdata <= 8'h00;
			14'd92: ff_rdata <= 8'h00;
			14'd93: ff_rdata <= 8'h00;
			14'd94: ff_rdata <= 8'h00;
			14'd95: ff_rdata <= 8'h00;
			14'd96: ff_rdata <= 8'h00;
			14'd97: ff_rdata <= 8'h00;
			14'd98: ff_rdata <= 8'h00;
			14'd99: ff_rdata <= 8'h00;
			14'd100: ff_rdata <= 8'h00;
			14'd101: ff_rdata <= 8'h00;
			14'd102: ff_rdata <= 8'h00;
			14'd103: ff_rdata <= 8'h00;
			14'd104: ff_rdata <= 8'h00;
			14'd105: ff_rdata <= 8'h00;
			14'd106: ff_rdata <= 8'h00;
			14'd107: ff_rdata <= 8'h00;
			14'd108: ff_rdata <= 8'h00;
			14'd109: ff_rdata <= 8'h00;
			14'd110: ff_rdata <= 8'h00;
			14'd111: ff_rdata <= 8'h00;
			14'd112: ff_rdata <= 8'h00;
			14'd113: ff_rdata <= 8'h00;
			14'd114: ff_rdata <= 8'h00;
			14'd115: ff_rdata <= 8'h00;
			14'd116: ff_rdata <= 8'h00;
			14'd117: ff_rdata <= 8'h00;
			14'd118: ff_rdata <= 8'h00;
			14'd119: ff_rdata <= 8'h00;
			14'd120: ff_rdata <= 8'h00;
			14'd121: ff_rdata <= 8'h00;
			14'd122: ff_rdata <= 8'h00;
			14'd123: ff_rdata <= 8'h00;
			14'd124: ff_rdata <= 8'h00;
			14'd125: ff_rdata <= 8'h00;
			14'd126: ff_rdata <= 8'h00;
			14'd127: ff_rdata <= 8'h00;
			14'd128: ff_rdata <= 8'h00;
			14'd129: ff_rdata <= 8'h00;
			14'd130: ff_rdata <= 8'h00;
			14'd131: ff_rdata <= 8'h00;
			14'd132: ff_rdata <= 8'h00;
			14'd133: ff_rdata <= 8'h00;
			14'd134: ff_rdata <= 8'h00;
			14'd135: ff_rdata <= 8'h00;
			14'd136: ff_rdata <= 8'h00;
			14'd137: ff_rdata <= 8'h00;
			14'd138: ff_rdata <= 8'h00;
			14'd139: ff_rdata <= 8'h00;
			14'd140: ff_rdata <= 8'h00;
			14'd141: ff_rdata <= 8'h00;
			14'd142: ff_rdata <= 8'h00;
			14'd143: ff_rdata <= 8'h00;
			14'd144: ff_rdata <= 8'h00;
			14'd145: ff_rdata <= 8'h00;
			14'd146: ff_rdata <= 8'h00;
			14'd147: ff_rdata <= 8'h00;
			14'd148: ff_rdata <= 8'h00;
			14'd149: ff_rdata <= 8'h00;
			14'd150: ff_rdata <= 8'h00;
			14'd151: ff_rdata <= 8'h00;
			14'd152: ff_rdata <= 8'h00;
			14'd153: ff_rdata <= 8'h00;
			14'd154: ff_rdata <= 8'h00;
			14'd155: ff_rdata <= 8'h00;
			14'd156: ff_rdata <= 8'h00;
			14'd157: ff_rdata <= 8'h00;
			14'd158: ff_rdata <= 8'h00;
			14'd159: ff_rdata <= 8'h00;
			14'd160: ff_rdata <= 8'h00;
			14'd161: ff_rdata <= 8'h00;
			14'd162: ff_rdata <= 8'h00;
			14'd163: ff_rdata <= 8'h00;
			14'd164: ff_rdata <= 8'h00;
			14'd165: ff_rdata <= 8'h00;
			14'd166: ff_rdata <= 8'h00;
			14'd167: ff_rdata <= 8'h00;
			14'd168: ff_rdata <= 8'h00;
			14'd169: ff_rdata <= 8'h00;
			14'd170: ff_rdata <= 8'h00;
			14'd171: ff_rdata <= 8'h00;
			14'd172: ff_rdata <= 8'h00;
			14'd173: ff_rdata <= 8'h00;
			14'd174: ff_rdata <= 8'h00;
			14'd175: ff_rdata <= 8'h00;
			14'd176: ff_rdata <= 8'h00;
			14'd177: ff_rdata <= 8'h00;
			14'd178: ff_rdata <= 8'h00;
			14'd179: ff_rdata <= 8'h00;
			14'd180: ff_rdata <= 8'h00;
			14'd181: ff_rdata <= 8'h00;
			14'd182: ff_rdata <= 8'h00;
			14'd183: ff_rdata <= 8'h00;
			14'd184: ff_rdata <= 8'h00;
			14'd185: ff_rdata <= 8'h00;
			14'd186: ff_rdata <= 8'h00;
			14'd187: ff_rdata <= 8'h00;
			14'd188: ff_rdata <= 8'h00;
			14'd189: ff_rdata <= 8'h00;
			14'd190: ff_rdata <= 8'h00;
			14'd191: ff_rdata <= 8'h00;
			14'd192: ff_rdata <= 8'h00;
			14'd193: ff_rdata <= 8'h00;
			14'd194: ff_rdata <= 8'h00;
			14'd195: ff_rdata <= 8'h00;
			14'd196: ff_rdata <= 8'h00;
			14'd197: ff_rdata <= 8'h00;
			14'd198: ff_rdata <= 8'h00;
			14'd199: ff_rdata <= 8'h00;
			14'd200: ff_rdata <= 8'h00;
			14'd201: ff_rdata <= 8'h00;
			14'd202: ff_rdata <= 8'h00;
			14'd203: ff_rdata <= 8'h00;
			14'd204: ff_rdata <= 8'h00;
			14'd205: ff_rdata <= 8'h00;
			14'd206: ff_rdata <= 8'h00;
			14'd207: ff_rdata <= 8'h00;
			14'd208: ff_rdata <= 8'h00;
			14'd209: ff_rdata <= 8'h00;
			14'd210: ff_rdata <= 8'h00;
			14'd211: ff_rdata <= 8'h00;
			14'd212: ff_rdata <= 8'h00;
			14'd213: ff_rdata <= 8'h00;
			14'd214: ff_rdata <= 8'h00;
			14'd215: ff_rdata <= 8'h00;
			14'd216: ff_rdata <= 8'h00;
			14'd217: ff_rdata <= 8'h00;
			14'd218: ff_rdata <= 8'h00;
			14'd219: ff_rdata <= 8'h00;
			14'd220: ff_rdata <= 8'h00;
			14'd221: ff_rdata <= 8'h00;
			14'd222: ff_rdata <= 8'h00;
			14'd223: ff_rdata <= 8'h00;
			14'd224: ff_rdata <= 8'h00;
			14'd225: ff_rdata <= 8'h00;
			14'd226: ff_rdata <= 8'h00;
			14'd227: ff_rdata <= 8'h00;
			14'd228: ff_rdata <= 8'h00;
			14'd229: ff_rdata <= 8'h00;
			14'd230: ff_rdata <= 8'h00;
			14'd231: ff_rdata <= 8'h00;
			14'd232: ff_rdata <= 8'h00;
			14'd233: ff_rdata <= 8'h00;
			14'd234: ff_rdata <= 8'h00;
			14'd235: ff_rdata <= 8'h00;
			14'd236: ff_rdata <= 8'h00;
			14'd237: ff_rdata <= 8'h00;
			14'd238: ff_rdata <= 8'h00;
			14'd239: ff_rdata <= 8'h00;
			14'd240: ff_rdata <= 8'h00;
			14'd241: ff_rdata <= 8'h00;
			14'd242: ff_rdata <= 8'h00;
			14'd243: ff_rdata <= 8'h00;
			14'd244: ff_rdata <= 8'h00;
			14'd245: ff_rdata <= 8'h00;
			14'd246: ff_rdata <= 8'h00;
			14'd247: ff_rdata <= 8'h00;
			14'd248: ff_rdata <= 8'h00;
			14'd249: ff_rdata <= 8'h00;
			14'd250: ff_rdata <= 8'h00;
			14'd251: ff_rdata <= 8'h00;
			14'd252: ff_rdata <= 8'h00;
			14'd253: ff_rdata <= 8'h00;
			14'd254: ff_rdata <= 8'h00;
			14'd255: ff_rdata <= 8'h00;
			14'd256: ff_rdata <= 8'h31;
			14'd257: ff_rdata <= 8'h00;
			14'd258: ff_rdata <= 8'h80;
			14'd259: ff_rdata <= 8'h21;
			14'd260: ff_rdata <= 8'hCC;
			14'd261: ff_rdata <= 8'h01;
			14'd262: ff_rdata <= 8'hCD;
			14'd263: ff_rdata <= 8'h8F;
			14'd264: ff_rdata <= 8'h01;
			14'd265: ff_rdata <= 8'h21;
			14'd266: ff_rdata <= 8'hD9;
			14'd267: ff_rdata <= 8'h01;
			14'd268: ff_rdata <= 8'hCD;
			14'd269: ff_rdata <= 8'h8F;
			14'd270: ff_rdata <= 8'h01;
			14'd271: ff_rdata <= 8'h01;
			14'd272: ff_rdata <= 8'h00;
			14'd273: ff_rdata <= 8'h00;
			14'd274: ff_rdata <= 8'hCD;
			14'd275: ff_rdata <= 8'h98;
			14'd276: ff_rdata <= 8'h01;
			14'd277: ff_rdata <= 8'h01;
			14'd278: ff_rdata <= 8'h01;
			14'd279: ff_rdata <= 8'h63;
			14'd280: ff_rdata <= 8'hCD;
			14'd281: ff_rdata <= 8'h98;
			14'd282: ff_rdata <= 8'h01;
			14'd283: ff_rdata <= 8'h01;
			14'd284: ff_rdata <= 8'h02;
			14'd285: ff_rdata <= 8'h06;
			14'd286: ff_rdata <= 8'hCD;
			14'd287: ff_rdata <= 8'h98;
			14'd288: ff_rdata <= 8'h01;
			14'd289: ff_rdata <= 8'h01;
			14'd290: ff_rdata <= 8'h03;
			14'd291: ff_rdata <= 8'h80;
			14'd292: ff_rdata <= 8'hCD;
			14'd293: ff_rdata <= 8'h98;
			14'd294: ff_rdata <= 8'h01;
			14'd295: ff_rdata <= 8'h01;
			14'd296: ff_rdata <= 8'h04;
			14'd297: ff_rdata <= 8'h00;
			14'd298: ff_rdata <= 8'hCD;
			14'd299: ff_rdata <= 8'h98;
			14'd300: ff_rdata <= 8'h01;
			14'd301: ff_rdata <= 8'h01;
			14'd302: ff_rdata <= 8'h05;
			14'd303: ff_rdata <= 8'h36;
			14'd304: ff_rdata <= 8'hCD;
			14'd305: ff_rdata <= 8'h98;
			14'd306: ff_rdata <= 8'h01;
			14'd307: ff_rdata <= 8'h01;
			14'd308: ff_rdata <= 8'h06;
			14'd309: ff_rdata <= 8'h07;
			14'd310: ff_rdata <= 8'hCD;
			14'd311: ff_rdata <= 8'h98;
			14'd312: ff_rdata <= 8'h01;
			14'd313: ff_rdata <= 8'h01;
			14'd314: ff_rdata <= 8'h07;
			14'd315: ff_rdata <= 8'hF7;
			14'd316: ff_rdata <= 8'hCD;
			14'd317: ff_rdata <= 8'h98;
			14'd318: ff_rdata <= 8'h01;
			14'd319: ff_rdata <= 8'h21;
			14'd320: ff_rdata <= 8'hEA;
			14'd321: ff_rdata <= 8'h01;
			14'd322: ff_rdata <= 8'hCD;
			14'd323: ff_rdata <= 8'h8F;
			14'd324: ff_rdata <= 8'h01;
			14'd325: ff_rdata <= 8'h21;
			14'd326: ff_rdata <= 8'h01;
			14'd327: ff_rdata <= 8'h02;
			14'd328: ff_rdata <= 8'hCD;
			14'd329: ff_rdata <= 8'h8F;
			14'd330: ff_rdata <= 8'h01;
			14'd331: ff_rdata <= 8'h21;
			14'd332: ff_rdata <= 8'h00;
			14'd333: ff_rdata <= 8'h00;
			14'd334: ff_rdata <= 8'h01;
			14'd335: ff_rdata <= 8'h00;
			14'd336: ff_rdata <= 8'h40;
			14'd337: ff_rdata <= 8'hAF;
			14'd338: ff_rdata <= 8'hCD;
			14'd339: ff_rdata <= 8'hAC;
			14'd340: ff_rdata <= 8'h01;
			14'd341: ff_rdata <= 8'h21;
			14'd342: ff_rdata <= 8'h00;
			14'd343: ff_rdata <= 8'h20;
			14'd344: ff_rdata <= 8'h01;
			14'd345: ff_rdata <= 8'h20;
			14'd346: ff_rdata <= 8'h00;
			14'd347: ff_rdata <= 8'h3E;
			14'd348: ff_rdata <= 8'hF4;
			14'd349: ff_rdata <= 8'hCD;
			14'd350: ff_rdata <= 8'hAC;
			14'd351: ff_rdata <= 8'h01;
			14'd352: ff_rdata <= 8'h21;
			14'd353: ff_rdata <= 8'hFE;
			14'd354: ff_rdata <= 8'h02;
			14'd355: ff_rdata <= 8'h11;
			14'd356: ff_rdata <= 8'h00;
			14'd357: ff_rdata <= 8'h00;
			14'd358: ff_rdata <= 8'h01;
			14'd359: ff_rdata <= 8'h00;
			14'd360: ff_rdata <= 8'h08;
			14'd361: ff_rdata <= 8'hCD;
			14'd362: ff_rdata <= 8'hBD;
			14'd363: ff_rdata <= 8'h01;
			14'd364: ff_rdata <= 8'h21;
			14'd365: ff_rdata <= 8'h1B;
			14'd366: ff_rdata <= 8'h02;
			14'd367: ff_rdata <= 8'h11;
			14'd368: ff_rdata <= 8'h00;
			14'd369: ff_rdata <= 8'h18;
			14'd370: ff_rdata <= 8'h01;
			14'd371: ff_rdata <= 8'hE3;
			14'd372: ff_rdata <= 8'h00;
			14'd373: ff_rdata <= 8'hCD;
			14'd374: ff_rdata <= 8'hBD;
			14'd375: ff_rdata <= 8'h01;
			14'd376: ff_rdata <= 8'h21;
			14'd377: ff_rdata <= 8'h11;
			14'd378: ff_rdata <= 8'h02;
			14'd379: ff_rdata <= 8'hCD;
			14'd380: ff_rdata <= 8'h8F;
			14'd381: ff_rdata <= 8'h01;
			14'd382: ff_rdata <= 8'h76;
			14'd383: ff_rdata <= 8'hDB;
			14'd384: ff_rdata <= 8'h10;
			14'd385: ff_rdata <= 8'h07;
			14'd386: ff_rdata <= 8'h07;
			14'd387: ff_rdata <= 8'hC9;
			14'd388: ff_rdata <= 8'h0E;
			14'd389: ff_rdata <= 8'h10;
			14'd390: ff_rdata <= 8'hED;
			14'd391: ff_rdata <= 8'h40;
			14'd392: ff_rdata <= 8'hCB;
			14'd393: ff_rdata <= 8'h18;
			14'd394: ff_rdata <= 8'h38;
			14'd395: ff_rdata <= 8'hFA;
			14'd396: ff_rdata <= 8'hED;
			14'd397: ff_rdata <= 8'h79;
			14'd398: ff_rdata <= 8'hC9;
			14'd399: ff_rdata <= 8'h7E;
			14'd400: ff_rdata <= 8'h23;
			14'd401: ff_rdata <= 8'hB7;
			14'd402: ff_rdata <= 8'hC8;
			14'd403: ff_rdata <= 8'hCD;
			14'd404: ff_rdata <= 8'h84;
			14'd405: ff_rdata <= 8'h01;
			14'd406: ff_rdata <= 8'h18;
			14'd407: ff_rdata <= 8'hF7;
			14'd408: ff_rdata <= 8'h78;
			14'd409: ff_rdata <= 8'hD3;
			14'd410: ff_rdata <= 8'h99;
			14'd411: ff_rdata <= 8'h79;
			14'd412: ff_rdata <= 8'hF6;
			14'd413: ff_rdata <= 8'h80;
			14'd414: ff_rdata <= 8'hD3;
			14'd415: ff_rdata <= 8'h99;
			14'd416: ff_rdata <= 8'hC9;
			14'd417: ff_rdata <= 8'h7D;
			14'd418: ff_rdata <= 8'hD3;
			14'd419: ff_rdata <= 8'h99;
			14'd420: ff_rdata <= 8'h7C;
			14'd421: ff_rdata <= 8'hE6;
			14'd422: ff_rdata <= 8'h3F;
			14'd423: ff_rdata <= 8'hF6;
			14'd424: ff_rdata <= 8'h40;
			14'd425: ff_rdata <= 8'hD3;
			14'd426: ff_rdata <= 8'h99;
			14'd427: ff_rdata <= 8'hC9;
			14'd428: ff_rdata <= 8'hF5;
			14'd429: ff_rdata <= 8'hCD;
			14'd430: ff_rdata <= 8'hA1;
			14'd431: ff_rdata <= 8'h01;
			14'd432: ff_rdata <= 8'hF1;
			14'd433: ff_rdata <= 8'hE5;
			14'd434: ff_rdata <= 8'h6F;
			14'd435: ff_rdata <= 8'h7D;
			14'd436: ff_rdata <= 8'hD3;
			14'd437: ff_rdata <= 8'h98;
			14'd438: ff_rdata <= 8'h0B;
			14'd439: ff_rdata <= 8'h79;
			14'd440: ff_rdata <= 8'hB0;
			14'd441: ff_rdata <= 8'h20;
			14'd442: ff_rdata <= 8'hF8;
			14'd443: ff_rdata <= 8'hE1;
			14'd444: ff_rdata <= 8'hC9;
			14'd445: ff_rdata <= 8'hEB;
			14'd446: ff_rdata <= 8'hCD;
			14'd447: ff_rdata <= 8'hA1;
			14'd448: ff_rdata <= 8'h01;
			14'd449: ff_rdata <= 8'hEB;
			14'd450: ff_rdata <= 8'h7E;
			14'd451: ff_rdata <= 8'h23;
			14'd452: ff_rdata <= 8'hD3;
			14'd453: ff_rdata <= 8'h98;
			14'd454: ff_rdata <= 8'h0B;
			14'd455: ff_rdata <= 8'h79;
			14'd456: ff_rdata <= 8'hB0;
			14'd457: ff_rdata <= 8'h20;
			14'd458: ff_rdata <= 8'hF7;
			14'd459: ff_rdata <= 8'hC9;
			14'd460: ff_rdata <= 8'h53;
			14'd461: ff_rdata <= 8'h74;
			14'd462: ff_rdata <= 8'h61;
			14'd463: ff_rdata <= 8'h72;
			14'd464: ff_rdata <= 8'h74;
			14'd465: ff_rdata <= 8'h20;
			14'd466: ff_rdata <= 8'h44;
			14'd467: ff_rdata <= 8'h45;
			14'd468: ff_rdata <= 8'h4D;
			14'd469: ff_rdata <= 8'h4F;
			14'd470: ff_rdata <= 8'h0D;
			14'd471: ff_rdata <= 8'h0A;
			14'd472: ff_rdata <= 8'h00;
			14'd473: ff_rdata <= 8'h2D;
			14'd474: ff_rdata <= 8'h2D;
			14'd475: ff_rdata <= 8'h20;
			14'd476: ff_rdata <= 8'h73;
			14'd477: ff_rdata <= 8'h65;
			14'd478: ff_rdata <= 8'h74;
			14'd479: ff_rdata <= 8'h20;
			14'd480: ff_rdata <= 8'h53;
			14'd481: ff_rdata <= 8'h43;
			14'd482: ff_rdata <= 8'h52;
			14'd483: ff_rdata <= 8'h45;
			14'd484: ff_rdata <= 8'h45;
			14'd485: ff_rdata <= 8'h4E;
			14'd486: ff_rdata <= 8'h31;
			14'd487: ff_rdata <= 8'h0D;
			14'd488: ff_rdata <= 8'h0A;
			14'd489: ff_rdata <= 8'h00;
			14'd490: ff_rdata <= 8'h2D;
			14'd491: ff_rdata <= 8'h2D;
			14'd492: ff_rdata <= 8'h20;
			14'd493: ff_rdata <= 8'h73;
			14'd494: ff_rdata <= 8'h65;
			14'd495: ff_rdata <= 8'h74;
			14'd496: ff_rdata <= 8'h20;
			14'd497: ff_rdata <= 8'h43;
			14'd498: ff_rdata <= 8'h4F;
			14'd499: ff_rdata <= 8'h4C;
			14'd500: ff_rdata <= 8'h4F;
			14'd501: ff_rdata <= 8'h52;
			14'd502: ff_rdata <= 8'h20;
			14'd503: ff_rdata <= 8'h50;
			14'd504: ff_rdata <= 8'h41;
			14'd505: ff_rdata <= 8'h4C;
			14'd506: ff_rdata <= 8'h45;
			14'd507: ff_rdata <= 8'h54;
			14'd508: ff_rdata <= 8'h54;
			14'd509: ff_rdata <= 8'h45;
			14'd510: ff_rdata <= 8'h0D;
			14'd511: ff_rdata <= 8'h0A;
			14'd512: ff_rdata <= 8'h00;
			14'd513: ff_rdata <= 8'h2D;
			14'd514: ff_rdata <= 8'h2D;
			14'd515: ff_rdata <= 8'h20;
			14'd516: ff_rdata <= 8'h63;
			14'd517: ff_rdata <= 8'h6C;
			14'd518: ff_rdata <= 8'h65;
			14'd519: ff_rdata <= 8'h61;
			14'd520: ff_rdata <= 8'h72;
			14'd521: ff_rdata <= 8'h20;
			14'd522: ff_rdata <= 8'h56;
			14'd523: ff_rdata <= 8'h52;
			14'd524: ff_rdata <= 8'h41;
			14'd525: ff_rdata <= 8'h4D;
			14'd526: ff_rdata <= 8'h0D;
			14'd527: ff_rdata <= 8'h0A;
			14'd528: ff_rdata <= 8'h00;
			14'd529: ff_rdata <= 8'h46;
			14'd530: ff_rdata <= 8'h69;
			14'd531: ff_rdata <= 8'h6E;
			14'd532: ff_rdata <= 8'h69;
			14'd533: ff_rdata <= 8'h73;
			14'd534: ff_rdata <= 8'h68;
			14'd535: ff_rdata <= 8'h2E;
			14'd536: ff_rdata <= 8'h0D;
			14'd537: ff_rdata <= 8'h0A;
			14'd538: ff_rdata <= 8'h00;
			14'd539: ff_rdata <= 8'h20;
			14'd540: ff_rdata <= 8'h20;
			14'd541: ff_rdata <= 8'h4D;
			14'd542: ff_rdata <= 8'h53;
			14'd543: ff_rdata <= 8'h58;
			14'd544: ff_rdata <= 8'h2D;
			14'd545: ff_rdata <= 8'h42;
			14'd546: ff_rdata <= 8'h41;
			14'd547: ff_rdata <= 8'h53;
			14'd548: ff_rdata <= 8'h49;
			14'd549: ff_rdata <= 8'h43;
			14'd550: ff_rdata <= 8'h20;
			14'd551: ff_rdata <= 8'h76;
			14'd552: ff_rdata <= 8'h65;
			14'd553: ff_rdata <= 8'h72;
			14'd554: ff_rdata <= 8'h73;
			14'd555: ff_rdata <= 8'h69;
			14'd556: ff_rdata <= 8'h6F;
			14'd557: ff_rdata <= 8'h6E;
			14'd558: ff_rdata <= 8'h20;
			14'd559: ff_rdata <= 8'h35;
			14'd560: ff_rdata <= 8'h2E;
			14'd561: ff_rdata <= 8'h30;
			14'd562: ff_rdata <= 8'h20;
			14'd563: ff_rdata <= 8'h20;
			14'd564: ff_rdata <= 8'h20;
			14'd565: ff_rdata <= 8'h20;
			14'd566: ff_rdata <= 8'h20;
			14'd567: ff_rdata <= 8'h20;
			14'd568: ff_rdata <= 8'h20;
			14'd569: ff_rdata <= 8'h20;
			14'd570: ff_rdata <= 8'h20;
			14'd571: ff_rdata <= 8'h20;
			14'd572: ff_rdata <= 8'h20;
			14'd573: ff_rdata <= 8'h43;
			14'd574: ff_rdata <= 8'h6F;
			14'd575: ff_rdata <= 8'h70;
			14'd576: ff_rdata <= 8'h79;
			14'd577: ff_rdata <= 8'h72;
			14'd578: ff_rdata <= 8'h69;
			14'd579: ff_rdata <= 8'h67;
			14'd580: ff_rdata <= 8'h68;
			14'd581: ff_rdata <= 8'h74;
			14'd582: ff_rdata <= 8'h20;
			14'd583: ff_rdata <= 8'h32;
			14'd584: ff_rdata <= 8'h30;
			14'd585: ff_rdata <= 8'h32;
			14'd586: ff_rdata <= 8'h35;
			14'd587: ff_rdata <= 8'h20;
			14'd588: ff_rdata <= 8'h62;
			14'd589: ff_rdata <= 8'h79;
			14'd590: ff_rdata <= 8'h20;
			14'd591: ff_rdata <= 8'h4D;
			14'd592: ff_rdata <= 8'h69;
			14'd593: ff_rdata <= 8'h63;
			14'd594: ff_rdata <= 8'h72;
			14'd595: ff_rdata <= 8'h6F;
			14'd596: ff_rdata <= 8'h73;
			14'd597: ff_rdata <= 8'h6F;
			14'd598: ff_rdata <= 8'h66;
			14'd599: ff_rdata <= 8'h74;
			14'd600: ff_rdata <= 8'h20;
			14'd601: ff_rdata <= 8'h20;
			14'd602: ff_rdata <= 8'h20;
			14'd603: ff_rdata <= 8'h20;
			14'd604: ff_rdata <= 8'h20;
			14'd605: ff_rdata <= 8'h49;
			14'd606: ff_rdata <= 8'h6F;
			14'd607: ff_rdata <= 8'h54;
			14'd608: ff_rdata <= 8'h20;
			14'd609: ff_rdata <= 8'h4D;
			14'd610: ff_rdata <= 8'h65;
			14'd611: ff_rdata <= 8'h64;
			14'd612: ff_rdata <= 8'h69;
			14'd613: ff_rdata <= 8'h61;
			14'd614: ff_rdata <= 8'h20;
			14'd615: ff_rdata <= 8'h4C;
			14'd616: ff_rdata <= 8'h61;
			14'd617: ff_rdata <= 8'h62;
			14'd618: ff_rdata <= 8'h20;
			14'd619: ff_rdata <= 8'h32;
			14'd620: ff_rdata <= 8'h30;
			14'd621: ff_rdata <= 8'h32;
			14'd622: ff_rdata <= 8'h35;
			14'd623: ff_rdata <= 8'h20;
			14'd624: ff_rdata <= 8'h20;
			14'd625: ff_rdata <= 8'h20;
			14'd626: ff_rdata <= 8'h20;
			14'd627: ff_rdata <= 8'h20;
			14'd628: ff_rdata <= 8'h20;
			14'd629: ff_rdata <= 8'h20;
			14'd630: ff_rdata <= 8'h20;
			14'd631: ff_rdata <= 8'h20;
			14'd632: ff_rdata <= 8'h20;
			14'd633: ff_rdata <= 8'h20;
			14'd634: ff_rdata <= 8'h20;
			14'd635: ff_rdata <= 8'h20;
			14'd636: ff_rdata <= 8'h20;
			14'd637: ff_rdata <= 8'h4D;
			14'd638: ff_rdata <= 8'h53;
			14'd639: ff_rdata <= 8'h58;
			14'd640: ff_rdata <= 8'h20;
			14'd641: ff_rdata <= 8'h4C;
			14'd642: ff_rdata <= 8'h69;
			14'd643: ff_rdata <= 8'h63;
			14'd644: ff_rdata <= 8'h65;
			14'd645: ff_rdata <= 8'h6E;
			14'd646: ff_rdata <= 8'h73;
			14'd647: ff_rdata <= 8'h69;
			14'd648: ff_rdata <= 8'h6E;
			14'd649: ff_rdata <= 8'h67;
			14'd650: ff_rdata <= 8'h20;
			14'd651: ff_rdata <= 8'h43;
			14'd652: ff_rdata <= 8'h6F;
			14'd653: ff_rdata <= 8'h72;
			14'd654: ff_rdata <= 8'h70;
			14'd655: ff_rdata <= 8'h20;
			14'd656: ff_rdata <= 8'h32;
			14'd657: ff_rdata <= 8'h30;
			14'd658: ff_rdata <= 8'h32;
			14'd659: ff_rdata <= 8'h35;
			14'd660: ff_rdata <= 8'h20;
			14'd661: ff_rdata <= 8'h20;
			14'd662: ff_rdata <= 8'h20;
			14'd663: ff_rdata <= 8'h20;
			14'd664: ff_rdata <= 8'h20;
			14'd665: ff_rdata <= 8'h20;
			14'd666: ff_rdata <= 8'h20;
			14'd667: ff_rdata <= 8'h20;
			14'd668: ff_rdata <= 8'h20;
			14'd669: ff_rdata <= 8'h32;
			14'd670: ff_rdata <= 8'h35;
			14'd671: ff_rdata <= 8'h32;
			14'd672: ff_rdata <= 8'h37;
			14'd673: ff_rdata <= 8'h31;
			14'd674: ff_rdata <= 8'h20;
			14'd675: ff_rdata <= 8'h42;
			14'd676: ff_rdata <= 8'h79;
			14'd677: ff_rdata <= 8'h74;
			14'd678: ff_rdata <= 8'h65;
			14'd679: ff_rdata <= 8'h73;
			14'd680: ff_rdata <= 8'h20;
			14'd681: ff_rdata <= 8'h66;
			14'd682: ff_rdata <= 8'h72;
			14'd683: ff_rdata <= 8'h65;
			14'd684: ff_rdata <= 8'h65;
			14'd685: ff_rdata <= 8'h20;
			14'd686: ff_rdata <= 8'h20;
			14'd687: ff_rdata <= 8'h20;
			14'd688: ff_rdata <= 8'h20;
			14'd689: ff_rdata <= 8'h20;
			14'd690: ff_rdata <= 8'h20;
			14'd691: ff_rdata <= 8'h20;
			14'd692: ff_rdata <= 8'h20;
			14'd693: ff_rdata <= 8'h20;
			14'd694: ff_rdata <= 8'h20;
			14'd695: ff_rdata <= 8'h20;
			14'd696: ff_rdata <= 8'h20;
			14'd697: ff_rdata <= 8'h20;
			14'd698: ff_rdata <= 8'h20;
			14'd699: ff_rdata <= 8'h20;
			14'd700: ff_rdata <= 8'h20;
			14'd701: ff_rdata <= 8'h44;
			14'd702: ff_rdata <= 8'h69;
			14'd703: ff_rdata <= 8'h73;
			14'd704: ff_rdata <= 8'h6B;
			14'd705: ff_rdata <= 8'h20;
			14'd706: ff_rdata <= 8'h42;
			14'd707: ff_rdata <= 8'h41;
			14'd708: ff_rdata <= 8'h53;
			14'd709: ff_rdata <= 8'h49;
			14'd710: ff_rdata <= 8'h43;
			14'd711: ff_rdata <= 8'h20;
			14'd712: ff_rdata <= 8'h76;
			14'd713: ff_rdata <= 8'h65;
			14'd714: ff_rdata <= 8'h72;
			14'd715: ff_rdata <= 8'h73;
			14'd716: ff_rdata <= 8'h69;
			14'd717: ff_rdata <= 8'h6F;
			14'd718: ff_rdata <= 8'h6E;
			14'd719: ff_rdata <= 8'h20;
			14'd720: ff_rdata <= 8'h33;
			14'd721: ff_rdata <= 8'h2E;
			14'd722: ff_rdata <= 8'h30;
			14'd723: ff_rdata <= 8'h30;
			14'd724: ff_rdata <= 8'h20;
			14'd725: ff_rdata <= 8'h20;
			14'd726: ff_rdata <= 8'h20;
			14'd727: ff_rdata <= 8'h20;
			14'd728: ff_rdata <= 8'h20;
			14'd729: ff_rdata <= 8'h20;
			14'd730: ff_rdata <= 8'h20;
			14'd731: ff_rdata <= 8'h20;
			14'd732: ff_rdata <= 8'h20;
			14'd733: ff_rdata <= 8'h4F;
			14'd734: ff_rdata <= 8'h6B;
			14'd735: ff_rdata <= 8'h20;
			14'd736: ff_rdata <= 8'h20;
			14'd737: ff_rdata <= 8'h20;
			14'd738: ff_rdata <= 8'h20;
			14'd739: ff_rdata <= 8'h20;
			14'd740: ff_rdata <= 8'h20;
			14'd741: ff_rdata <= 8'h20;
			14'd742: ff_rdata <= 8'h20;
			14'd743: ff_rdata <= 8'h20;
			14'd744: ff_rdata <= 8'h20;
			14'd745: ff_rdata <= 8'h20;
			14'd746: ff_rdata <= 8'h20;
			14'd747: ff_rdata <= 8'h20;
			14'd748: ff_rdata <= 8'h20;
			14'd749: ff_rdata <= 8'h20;
			14'd750: ff_rdata <= 8'h20;
			14'd751: ff_rdata <= 8'h20;
			14'd752: ff_rdata <= 8'h20;
			14'd753: ff_rdata <= 8'h20;
			14'd754: ff_rdata <= 8'h20;
			14'd755: ff_rdata <= 8'h20;
			14'd756: ff_rdata <= 8'h20;
			14'd757: ff_rdata <= 8'h20;
			14'd758: ff_rdata <= 8'h20;
			14'd759: ff_rdata <= 8'h20;
			14'd760: ff_rdata <= 8'h20;
			14'd761: ff_rdata <= 8'h20;
			14'd762: ff_rdata <= 8'h20;
			14'd763: ff_rdata <= 8'h20;
			14'd764: ff_rdata <= 8'h20;
			14'd765: ff_rdata <= 8'hFF;
			14'd766: ff_rdata <= 8'h00;
			14'd767: ff_rdata <= 8'h00;
			14'd768: ff_rdata <= 8'h00;
			14'd769: ff_rdata <= 8'h00;
			14'd770: ff_rdata <= 8'h00;
			14'd771: ff_rdata <= 8'h00;
			14'd772: ff_rdata <= 8'h00;
			14'd773: ff_rdata <= 8'h00;
			14'd774: ff_rdata <= 8'h7E;
			14'd775: ff_rdata <= 8'h42;
			14'd776: ff_rdata <= 8'h7E;
			14'd777: ff_rdata <= 8'h42;
			14'd778: ff_rdata <= 8'h7E;
			14'd779: ff_rdata <= 8'h42;
			14'd780: ff_rdata <= 8'h82;
			14'd781: ff_rdata <= 8'h00;
			14'd782: ff_rdata <= 8'h10;
			14'd783: ff_rdata <= 8'h92;
			14'd784: ff_rdata <= 8'h54;
			14'd785: ff_rdata <= 8'h10;
			14'd786: ff_rdata <= 8'h28;
			14'd787: ff_rdata <= 8'h44;
			14'd788: ff_rdata <= 8'h82;
			14'd789: ff_rdata <= 8'h00;
			14'd790: ff_rdata <= 8'h12;
			14'd791: ff_rdata <= 8'h14;
			14'd792: ff_rdata <= 8'hF8;
			14'd793: ff_rdata <= 8'h14;
			14'd794: ff_rdata <= 8'h34;
			14'd795: ff_rdata <= 8'h52;
			14'd796: ff_rdata <= 8'h92;
			14'd797: ff_rdata <= 8'h00;
			14'd798: ff_rdata <= 8'h10;
			14'd799: ff_rdata <= 8'h10;
			14'd800: ff_rdata <= 8'hFE;
			14'd801: ff_rdata <= 8'h10;
			14'd802: ff_rdata <= 8'h38;
			14'd803: ff_rdata <= 8'h54;
			14'd804: ff_rdata <= 8'h92;
			14'd805: ff_rdata <= 8'h00;
			14'd806: ff_rdata <= 8'h10;
			14'd807: ff_rdata <= 8'h28;
			14'd808: ff_rdata <= 8'h7C;
			14'd809: ff_rdata <= 8'h92;
			14'd810: ff_rdata <= 8'h38;
			14'd811: ff_rdata <= 8'h54;
			14'd812: ff_rdata <= 8'hFE;
			14'd813: ff_rdata <= 8'h00;
			14'd814: ff_rdata <= 8'h10;
			14'd815: ff_rdata <= 8'h10;
			14'd816: ff_rdata <= 8'h10;
			14'd817: ff_rdata <= 8'h7C;
			14'd818: ff_rdata <= 8'h10;
			14'd819: ff_rdata <= 8'h10;
			14'd820: ff_rdata <= 8'hFE;
			14'd821: ff_rdata <= 8'h00;
			14'd822: ff_rdata <= 8'h7E;
			14'd823: ff_rdata <= 8'h42;
			14'd824: ff_rdata <= 8'h42;
			14'd825: ff_rdata <= 8'h7E;
			14'd826: ff_rdata <= 8'h42;
			14'd827: ff_rdata <= 8'h42;
			14'd828: ff_rdata <= 8'h7E;
			14'd829: ff_rdata <= 8'h00;
			14'd830: ff_rdata <= 8'h40;
			14'd831: ff_rdata <= 8'h7E;
			14'd832: ff_rdata <= 8'h48;
			14'd833: ff_rdata <= 8'h3C;
			14'd834: ff_rdata <= 8'h28;
			14'd835: ff_rdata <= 8'h7E;
			14'd836: ff_rdata <= 8'h08;
			14'd837: ff_rdata <= 8'h00;
			14'd838: ff_rdata <= 8'hFE;
			14'd839: ff_rdata <= 8'h92;
			14'd840: ff_rdata <= 8'h92;
			14'd841: ff_rdata <= 8'hFE;
			14'd842: ff_rdata <= 8'h82;
			14'd843: ff_rdata <= 8'h82;
			14'd844: ff_rdata <= 8'h86;
			14'd845: ff_rdata <= 8'h00;
			14'd846: ff_rdata <= 8'h04;
			14'd847: ff_rdata <= 8'hEE;
			14'd848: ff_rdata <= 8'hA4;
			14'd849: ff_rdata <= 8'hEF;
			14'd850: ff_rdata <= 8'hA2;
			14'd851: ff_rdata <= 8'hEA;
			14'd852: ff_rdata <= 8'h06;
			14'd853: ff_rdata <= 8'h00;
			14'd854: ff_rdata <= 8'h28;
			14'd855: ff_rdata <= 8'h44;
			14'd856: ff_rdata <= 8'h82;
			14'd857: ff_rdata <= 8'h3C;
			14'd858: ff_rdata <= 8'h14;
			14'd859: ff_rdata <= 8'h24;
			14'd860: ff_rdata <= 8'h4C;
			14'd861: ff_rdata <= 8'h00;
			14'd862: ff_rdata <= 8'h28;
			14'd863: ff_rdata <= 8'hC8;
			14'd864: ff_rdata <= 8'h5C;
			14'd865: ff_rdata <= 8'hEA;
			14'd866: ff_rdata <= 8'h6C;
			14'd867: ff_rdata <= 8'hC8;
			14'd868: ff_rdata <= 8'h50;
			14'd869: ff_rdata <= 8'h00;
			14'd870: ff_rdata <= 8'h7C;
			14'd871: ff_rdata <= 8'h20;
			14'd872: ff_rdata <= 8'h7C;
			14'd873: ff_rdata <= 8'h44;
			14'd874: ff_rdata <= 8'h7C;
			14'd875: ff_rdata <= 8'h44;
			14'd876: ff_rdata <= 8'h7C;
			14'd877: ff_rdata <= 8'h00;
			14'd878: ff_rdata <= 8'h0C;
			14'd879: ff_rdata <= 8'h70;
			14'd880: ff_rdata <= 8'h10;
			14'd881: ff_rdata <= 8'hFE;
			14'd882: ff_rdata <= 8'h10;
			14'd883: ff_rdata <= 8'h10;
			14'd884: ff_rdata <= 8'h10;
			14'd885: ff_rdata <= 8'h00;
			14'd886: ff_rdata <= 8'h7E;
			14'd887: ff_rdata <= 8'h10;
			14'd888: ff_rdata <= 8'h1E;
			14'd889: ff_rdata <= 8'h12;
			14'd890: ff_rdata <= 8'h22;
			14'd891: ff_rdata <= 8'h44;
			14'd892: ff_rdata <= 8'h08;
			14'd893: ff_rdata <= 8'h00;
			14'd894: ff_rdata <= 8'h00;
			14'd895: ff_rdata <= 8'h7C;
			14'd896: ff_rdata <= 8'h28;
			14'd897: ff_rdata <= 8'h28;
			14'd898: ff_rdata <= 8'h28;
			14'd899: ff_rdata <= 8'h4E;
			14'd900: ff_rdata <= 8'h00;
			14'd901: ff_rdata <= 8'h00;
			14'd902: ff_rdata <= 8'h10;
			14'd903: ff_rdata <= 8'h10;
			14'd904: ff_rdata <= 8'h10;
			14'd905: ff_rdata <= 8'hFF;
			14'd906: ff_rdata <= 8'h00;
			14'd907: ff_rdata <= 8'h00;
			14'd908: ff_rdata <= 8'h00;
			14'd909: ff_rdata <= 8'h00;
			14'd910: ff_rdata <= 8'h00;
			14'd911: ff_rdata <= 8'h00;
			14'd912: ff_rdata <= 8'h00;
			14'd913: ff_rdata <= 8'hFF;
			14'd914: ff_rdata <= 8'h10;
			14'd915: ff_rdata <= 8'h10;
			14'd916: ff_rdata <= 8'h10;
			14'd917: ff_rdata <= 8'h10;
			14'd918: ff_rdata <= 8'h10;
			14'd919: ff_rdata <= 8'h10;
			14'd920: ff_rdata <= 8'h10;
			14'd921: ff_rdata <= 8'hF0;
			14'd922: ff_rdata <= 8'h10;
			14'd923: ff_rdata <= 8'h10;
			14'd924: ff_rdata <= 8'h10;
			14'd925: ff_rdata <= 8'h10;
			14'd926: ff_rdata <= 8'h10;
			14'd927: ff_rdata <= 8'h10;
			14'd928: ff_rdata <= 8'h10;
			14'd929: ff_rdata <= 8'h1F;
			14'd930: ff_rdata <= 8'h10;
			14'd931: ff_rdata <= 8'h10;
			14'd932: ff_rdata <= 8'h10;
			14'd933: ff_rdata <= 8'h10;
			14'd934: ff_rdata <= 8'h10;
			14'd935: ff_rdata <= 8'h10;
			14'd936: ff_rdata <= 8'h10;
			14'd937: ff_rdata <= 8'hFF;
			14'd938: ff_rdata <= 8'h10;
			14'd939: ff_rdata <= 8'h10;
			14'd940: ff_rdata <= 8'h10;
			14'd941: ff_rdata <= 8'h10;
			14'd942: ff_rdata <= 8'h10;
			14'd943: ff_rdata <= 8'h10;
			14'd944: ff_rdata <= 8'h10;
			14'd945: ff_rdata <= 8'h10;
			14'd946: ff_rdata <= 8'h10;
			14'd947: ff_rdata <= 8'h10;
			14'd948: ff_rdata <= 8'h10;
			14'd949: ff_rdata <= 8'h10;
			14'd950: ff_rdata <= 8'h00;
			14'd951: ff_rdata <= 8'h00;
			14'd952: ff_rdata <= 8'h00;
			14'd953: ff_rdata <= 8'hFF;
			14'd954: ff_rdata <= 8'h00;
			14'd955: ff_rdata <= 8'h00;
			14'd956: ff_rdata <= 8'h00;
			14'd957: ff_rdata <= 8'h00;
			14'd958: ff_rdata <= 8'h00;
			14'd959: ff_rdata <= 8'h00;
			14'd960: ff_rdata <= 8'h00;
			14'd961: ff_rdata <= 8'h1F;
			14'd962: ff_rdata <= 8'h10;
			14'd963: ff_rdata <= 8'h10;
			14'd964: ff_rdata <= 8'h10;
			14'd965: ff_rdata <= 8'h10;
			14'd966: ff_rdata <= 8'h00;
			14'd967: ff_rdata <= 8'h00;
			14'd968: ff_rdata <= 8'h00;
			14'd969: ff_rdata <= 8'hF0;
			14'd970: ff_rdata <= 8'h10;
			14'd971: ff_rdata <= 8'h10;
			14'd972: ff_rdata <= 8'h10;
			14'd973: ff_rdata <= 8'h10;
			14'd974: ff_rdata <= 8'h10;
			14'd975: ff_rdata <= 8'h10;
			14'd976: ff_rdata <= 8'h10;
			14'd977: ff_rdata <= 8'h1F;
			14'd978: ff_rdata <= 8'h00;
			14'd979: ff_rdata <= 8'h00;
			14'd980: ff_rdata <= 8'h00;
			14'd981: ff_rdata <= 8'h00;
			14'd982: ff_rdata <= 8'h10;
			14'd983: ff_rdata <= 8'h10;
			14'd984: ff_rdata <= 8'h10;
			14'd985: ff_rdata <= 8'hF0;
			14'd986: ff_rdata <= 8'h00;
			14'd987: ff_rdata <= 8'h00;
			14'd988: ff_rdata <= 8'h00;
			14'd989: ff_rdata <= 8'h00;
			14'd990: ff_rdata <= 8'h81;
			14'd991: ff_rdata <= 8'h42;
			14'd992: ff_rdata <= 8'h24;
			14'd993: ff_rdata <= 8'h18;
			14'd994: ff_rdata <= 8'h18;
			14'd995: ff_rdata <= 8'h24;
			14'd996: ff_rdata <= 8'h42;
			14'd997: ff_rdata <= 8'h81;
			14'd998: ff_rdata <= 8'h10;
			14'd999: ff_rdata <= 8'h7C;
			14'd1000: ff_rdata <= 8'h10;
			14'd1001: ff_rdata <= 8'h10;
			14'd1002: ff_rdata <= 8'h28;
			14'd1003: ff_rdata <= 8'h44;
			14'd1004: ff_rdata <= 8'h82;
			14'd1005: ff_rdata <= 8'h00;
			14'd1006: ff_rdata <= 8'h10;
			14'd1007: ff_rdata <= 8'h10;
			14'd1008: ff_rdata <= 8'hFE;
			14'd1009: ff_rdata <= 8'h92;
			14'd1010: ff_rdata <= 8'hFE;
			14'd1011: ff_rdata <= 8'h10;
			14'd1012: ff_rdata <= 8'h10;
			14'd1013: ff_rdata <= 8'h00;
			14'd1014: ff_rdata <= 8'h10;
			14'd1015: ff_rdata <= 8'h10;
			14'd1016: ff_rdata <= 8'h54;
			14'd1017: ff_rdata <= 8'h54;
			14'd1018: ff_rdata <= 8'h92;
			14'd1019: ff_rdata <= 8'h10;
			14'd1020: ff_rdata <= 8'h30;
			14'd1021: ff_rdata <= 8'h00;
			14'd1022: ff_rdata <= 8'h00;
			14'd1023: ff_rdata <= 8'h00;
			14'd1024: ff_rdata <= 8'h00;
			14'd1025: ff_rdata <= 8'h00;
			14'd1026: ff_rdata <= 8'h00;
			14'd1027: ff_rdata <= 8'h00;
			14'd1028: ff_rdata <= 8'h00;
			14'd1029: ff_rdata <= 8'h00;
			14'd1030: ff_rdata <= 8'h20;
			14'd1031: ff_rdata <= 8'h20;
			14'd1032: ff_rdata <= 8'h20;
			14'd1033: ff_rdata <= 8'h20;
			14'd1034: ff_rdata <= 8'h00;
			14'd1035: ff_rdata <= 8'h00;
			14'd1036: ff_rdata <= 8'h20;
			14'd1037: ff_rdata <= 8'h00;
			14'd1038: ff_rdata <= 8'h50;
			14'd1039: ff_rdata <= 8'h50;
			14'd1040: ff_rdata <= 8'h50;
			14'd1041: ff_rdata <= 8'h00;
			14'd1042: ff_rdata <= 8'h00;
			14'd1043: ff_rdata <= 8'h00;
			14'd1044: ff_rdata <= 8'h00;
			14'd1045: ff_rdata <= 8'h00;
			14'd1046: ff_rdata <= 8'h50;
			14'd1047: ff_rdata <= 8'h50;
			14'd1048: ff_rdata <= 8'hF8;
			14'd1049: ff_rdata <= 8'h50;
			14'd1050: ff_rdata <= 8'hF8;
			14'd1051: ff_rdata <= 8'h50;
			14'd1052: ff_rdata <= 8'h50;
			14'd1053: ff_rdata <= 8'h00;
			14'd1054: ff_rdata <= 8'h20;
			14'd1055: ff_rdata <= 8'h78;
			14'd1056: ff_rdata <= 8'hA0;
			14'd1057: ff_rdata <= 8'h70;
			14'd1058: ff_rdata <= 8'h28;
			14'd1059: ff_rdata <= 8'hF0;
			14'd1060: ff_rdata <= 8'h20;
			14'd1061: ff_rdata <= 8'h00;
			14'd1062: ff_rdata <= 8'hC0;
			14'd1063: ff_rdata <= 8'hC8;
			14'd1064: ff_rdata <= 8'h10;
			14'd1065: ff_rdata <= 8'h20;
			14'd1066: ff_rdata <= 8'h40;
			14'd1067: ff_rdata <= 8'h98;
			14'd1068: ff_rdata <= 8'h18;
			14'd1069: ff_rdata <= 8'h00;
			14'd1070: ff_rdata <= 8'h40;
			14'd1071: ff_rdata <= 8'hA0;
			14'd1072: ff_rdata <= 8'h40;
			14'd1073: ff_rdata <= 8'hA8;
			14'd1074: ff_rdata <= 8'h90;
			14'd1075: ff_rdata <= 8'h98;
			14'd1076: ff_rdata <= 8'h60;
			14'd1077: ff_rdata <= 8'h00;
			14'd1078: ff_rdata <= 8'h10;
			14'd1079: ff_rdata <= 8'h20;
			14'd1080: ff_rdata <= 8'h40;
			14'd1081: ff_rdata <= 8'h00;
			14'd1082: ff_rdata <= 8'h00;
			14'd1083: ff_rdata <= 8'h00;
			14'd1084: ff_rdata <= 8'h00;
			14'd1085: ff_rdata <= 8'h00;
			14'd1086: ff_rdata <= 8'h10;
			14'd1087: ff_rdata <= 8'h20;
			14'd1088: ff_rdata <= 8'h40;
			14'd1089: ff_rdata <= 8'h40;
			14'd1090: ff_rdata <= 8'h40;
			14'd1091: ff_rdata <= 8'h20;
			14'd1092: ff_rdata <= 8'h10;
			14'd1093: ff_rdata <= 8'h00;
			14'd1094: ff_rdata <= 8'h40;
			14'd1095: ff_rdata <= 8'h20;
			14'd1096: ff_rdata <= 8'h10;
			14'd1097: ff_rdata <= 8'h10;
			14'd1098: ff_rdata <= 8'h10;
			14'd1099: ff_rdata <= 8'h20;
			14'd1100: ff_rdata <= 8'h40;
			14'd1101: ff_rdata <= 8'h00;
			14'd1102: ff_rdata <= 8'h20;
			14'd1103: ff_rdata <= 8'hA8;
			14'd1104: ff_rdata <= 8'h70;
			14'd1105: ff_rdata <= 8'h20;
			14'd1106: ff_rdata <= 8'h70;
			14'd1107: ff_rdata <= 8'hA8;
			14'd1108: ff_rdata <= 8'h20;
			14'd1109: ff_rdata <= 8'h00;
			14'd1110: ff_rdata <= 8'h00;
			14'd1111: ff_rdata <= 8'h20;
			14'd1112: ff_rdata <= 8'h20;
			14'd1113: ff_rdata <= 8'hF8;
			14'd1114: ff_rdata <= 8'h20;
			14'd1115: ff_rdata <= 8'h20;
			14'd1116: ff_rdata <= 8'h00;
			14'd1117: ff_rdata <= 8'h00;
			14'd1118: ff_rdata <= 8'h00;
			14'd1119: ff_rdata <= 8'h00;
			14'd1120: ff_rdata <= 8'h00;
			14'd1121: ff_rdata <= 8'h00;
			14'd1122: ff_rdata <= 8'h00;
			14'd1123: ff_rdata <= 8'h20;
			14'd1124: ff_rdata <= 8'h20;
			14'd1125: ff_rdata <= 8'h40;
			14'd1126: ff_rdata <= 8'h00;
			14'd1127: ff_rdata <= 8'h00;
			14'd1128: ff_rdata <= 8'h00;
			14'd1129: ff_rdata <= 8'h78;
			14'd1130: ff_rdata <= 8'h00;
			14'd1131: ff_rdata <= 8'h00;
			14'd1132: ff_rdata <= 8'h00;
			14'd1133: ff_rdata <= 8'h00;
			14'd1134: ff_rdata <= 8'h00;
			14'd1135: ff_rdata <= 8'h00;
			14'd1136: ff_rdata <= 8'h00;
			14'd1137: ff_rdata <= 8'h00;
			14'd1138: ff_rdata <= 8'h00;
			14'd1139: ff_rdata <= 8'h60;
			14'd1140: ff_rdata <= 8'h60;
			14'd1141: ff_rdata <= 8'h00;
			14'd1142: ff_rdata <= 8'h00;
			14'd1143: ff_rdata <= 8'h00;
			14'd1144: ff_rdata <= 8'h08;
			14'd1145: ff_rdata <= 8'h10;
			14'd1146: ff_rdata <= 8'h20;
			14'd1147: ff_rdata <= 8'h40;
			14'd1148: ff_rdata <= 8'h80;
			14'd1149: ff_rdata <= 8'h00;
			14'd1150: ff_rdata <= 8'h70;
			14'd1151: ff_rdata <= 8'h88;
			14'd1152: ff_rdata <= 8'h98;
			14'd1153: ff_rdata <= 8'hA8;
			14'd1154: ff_rdata <= 8'hC8;
			14'd1155: ff_rdata <= 8'h88;
			14'd1156: ff_rdata <= 8'h70;
			14'd1157: ff_rdata <= 8'h00;
			14'd1158: ff_rdata <= 8'h20;
			14'd1159: ff_rdata <= 8'h60;
			14'd1160: ff_rdata <= 8'hA0;
			14'd1161: ff_rdata <= 8'h20;
			14'd1162: ff_rdata <= 8'h20;
			14'd1163: ff_rdata <= 8'h20;
			14'd1164: ff_rdata <= 8'hF8;
			14'd1165: ff_rdata <= 8'h00;
			14'd1166: ff_rdata <= 8'h70;
			14'd1167: ff_rdata <= 8'h88;
			14'd1168: ff_rdata <= 8'h08;
			14'd1169: ff_rdata <= 8'h10;
			14'd1170: ff_rdata <= 8'h60;
			14'd1171: ff_rdata <= 8'h80;
			14'd1172: ff_rdata <= 8'hF8;
			14'd1173: ff_rdata <= 8'h00;
			14'd1174: ff_rdata <= 8'h70;
			14'd1175: ff_rdata <= 8'h88;
			14'd1176: ff_rdata <= 8'h08;
			14'd1177: ff_rdata <= 8'h30;
			14'd1178: ff_rdata <= 8'h08;
			14'd1179: ff_rdata <= 8'h88;
			14'd1180: ff_rdata <= 8'h70;
			14'd1181: ff_rdata <= 8'h00;
			14'd1182: ff_rdata <= 8'h10;
			14'd1183: ff_rdata <= 8'h30;
			14'd1184: ff_rdata <= 8'h50;
			14'd1185: ff_rdata <= 8'h90;
			14'd1186: ff_rdata <= 8'hF8;
			14'd1187: ff_rdata <= 8'h10;
			14'd1188: ff_rdata <= 8'h10;
			14'd1189: ff_rdata <= 8'h00;
			14'd1190: ff_rdata <= 8'hF8;
			14'd1191: ff_rdata <= 8'h80;
			14'd1192: ff_rdata <= 8'hE0;
			14'd1193: ff_rdata <= 8'h10;
			14'd1194: ff_rdata <= 8'h08;
			14'd1195: ff_rdata <= 8'h10;
			14'd1196: ff_rdata <= 8'hE0;
			14'd1197: ff_rdata <= 8'h00;
			14'd1198: ff_rdata <= 8'h30;
			14'd1199: ff_rdata <= 8'h40;
			14'd1200: ff_rdata <= 8'h80;
			14'd1201: ff_rdata <= 8'hF0;
			14'd1202: ff_rdata <= 8'h88;
			14'd1203: ff_rdata <= 8'h88;
			14'd1204: ff_rdata <= 8'h70;
			14'd1205: ff_rdata <= 8'h00;
			14'd1206: ff_rdata <= 8'hF8;
			14'd1207: ff_rdata <= 8'h88;
			14'd1208: ff_rdata <= 8'h10;
			14'd1209: ff_rdata <= 8'h20;
			14'd1210: ff_rdata <= 8'h20;
			14'd1211: ff_rdata <= 8'h20;
			14'd1212: ff_rdata <= 8'h20;
			14'd1213: ff_rdata <= 8'h00;
			14'd1214: ff_rdata <= 8'h70;
			14'd1215: ff_rdata <= 8'h88;
			14'd1216: ff_rdata <= 8'h88;
			14'd1217: ff_rdata <= 8'h70;
			14'd1218: ff_rdata <= 8'h88;
			14'd1219: ff_rdata <= 8'h88;
			14'd1220: ff_rdata <= 8'h70;
			14'd1221: ff_rdata <= 8'h00;
			14'd1222: ff_rdata <= 8'h70;
			14'd1223: ff_rdata <= 8'h88;
			14'd1224: ff_rdata <= 8'h88;
			14'd1225: ff_rdata <= 8'h78;
			14'd1226: ff_rdata <= 8'h08;
			14'd1227: ff_rdata <= 8'h10;
			14'd1228: ff_rdata <= 8'h60;
			14'd1229: ff_rdata <= 8'h00;
			14'd1230: ff_rdata <= 8'h00;
			14'd1231: ff_rdata <= 8'h00;
			14'd1232: ff_rdata <= 8'h20;
			14'd1233: ff_rdata <= 8'h00;
			14'd1234: ff_rdata <= 8'h00;
			14'd1235: ff_rdata <= 8'h20;
			14'd1236: ff_rdata <= 8'h00;
			14'd1237: ff_rdata <= 8'h00;
			14'd1238: ff_rdata <= 8'h00;
			14'd1239: ff_rdata <= 8'h00;
			14'd1240: ff_rdata <= 8'h20;
			14'd1241: ff_rdata <= 8'h00;
			14'd1242: ff_rdata <= 8'h00;
			14'd1243: ff_rdata <= 8'h20;
			14'd1244: ff_rdata <= 8'h20;
			14'd1245: ff_rdata <= 8'h40;
			14'd1246: ff_rdata <= 8'h18;
			14'd1247: ff_rdata <= 8'h30;
			14'd1248: ff_rdata <= 8'h60;
			14'd1249: ff_rdata <= 8'hC0;
			14'd1250: ff_rdata <= 8'h60;
			14'd1251: ff_rdata <= 8'h30;
			14'd1252: ff_rdata <= 8'h18;
			14'd1253: ff_rdata <= 8'h00;
			14'd1254: ff_rdata <= 8'h00;
			14'd1255: ff_rdata <= 8'h00;
			14'd1256: ff_rdata <= 8'hF8;
			14'd1257: ff_rdata <= 8'h00;
			14'd1258: ff_rdata <= 8'hF8;
			14'd1259: ff_rdata <= 8'h00;
			14'd1260: ff_rdata <= 8'h00;
			14'd1261: ff_rdata <= 8'h00;
			14'd1262: ff_rdata <= 8'hC0;
			14'd1263: ff_rdata <= 8'h60;
			14'd1264: ff_rdata <= 8'h30;
			14'd1265: ff_rdata <= 8'h18;
			14'd1266: ff_rdata <= 8'h30;
			14'd1267: ff_rdata <= 8'h60;
			14'd1268: ff_rdata <= 8'hC0;
			14'd1269: ff_rdata <= 8'h00;
			14'd1270: ff_rdata <= 8'h70;
			14'd1271: ff_rdata <= 8'h88;
			14'd1272: ff_rdata <= 8'h08;
			14'd1273: ff_rdata <= 8'h10;
			14'd1274: ff_rdata <= 8'h20;
			14'd1275: ff_rdata <= 8'h00;
			14'd1276: ff_rdata <= 8'h20;
			14'd1277: ff_rdata <= 8'h00;
			14'd1278: ff_rdata <= 8'h70;
			14'd1279: ff_rdata <= 8'h88;
			14'd1280: ff_rdata <= 8'h08;
			14'd1281: ff_rdata <= 8'h68;
			14'd1282: ff_rdata <= 8'hA8;
			14'd1283: ff_rdata <= 8'hA8;
			14'd1284: ff_rdata <= 8'h70;
			14'd1285: ff_rdata <= 8'h00;
			14'd1286: ff_rdata <= 8'h20;
			14'd1287: ff_rdata <= 8'h50;
			14'd1288: ff_rdata <= 8'h88;
			14'd1289: ff_rdata <= 8'h88;
			14'd1290: ff_rdata <= 8'hF8;
			14'd1291: ff_rdata <= 8'h88;
			14'd1292: ff_rdata <= 8'h88;
			14'd1293: ff_rdata <= 8'h00;
			14'd1294: ff_rdata <= 8'hF0;
			14'd1295: ff_rdata <= 8'h48;
			14'd1296: ff_rdata <= 8'h48;
			14'd1297: ff_rdata <= 8'h70;
			14'd1298: ff_rdata <= 8'h48;
			14'd1299: ff_rdata <= 8'h48;
			14'd1300: ff_rdata <= 8'hF0;
			14'd1301: ff_rdata <= 8'h00;
			14'd1302: ff_rdata <= 8'h30;
			14'd1303: ff_rdata <= 8'h48;
			14'd1304: ff_rdata <= 8'h80;
			14'd1305: ff_rdata <= 8'h80;
			14'd1306: ff_rdata <= 8'h80;
			14'd1307: ff_rdata <= 8'h48;
			14'd1308: ff_rdata <= 8'h30;
			14'd1309: ff_rdata <= 8'h00;
			14'd1310: ff_rdata <= 8'hE0;
			14'd1311: ff_rdata <= 8'h50;
			14'd1312: ff_rdata <= 8'h48;
			14'd1313: ff_rdata <= 8'h48;
			14'd1314: ff_rdata <= 8'h48;
			14'd1315: ff_rdata <= 8'h50;
			14'd1316: ff_rdata <= 8'hE0;
			14'd1317: ff_rdata <= 8'h00;
			14'd1318: ff_rdata <= 8'hF8;
			14'd1319: ff_rdata <= 8'h80;
			14'd1320: ff_rdata <= 8'h80;
			14'd1321: ff_rdata <= 8'hF0;
			14'd1322: ff_rdata <= 8'h80;
			14'd1323: ff_rdata <= 8'h80;
			14'd1324: ff_rdata <= 8'hF8;
			14'd1325: ff_rdata <= 8'h00;
			14'd1326: ff_rdata <= 8'hF8;
			14'd1327: ff_rdata <= 8'h80;
			14'd1328: ff_rdata <= 8'h80;
			14'd1329: ff_rdata <= 8'hF0;
			14'd1330: ff_rdata <= 8'h80;
			14'd1331: ff_rdata <= 8'h80;
			14'd1332: ff_rdata <= 8'h80;
			14'd1333: ff_rdata <= 8'h00;
			14'd1334: ff_rdata <= 8'h70;
			14'd1335: ff_rdata <= 8'h88;
			14'd1336: ff_rdata <= 8'h80;
			14'd1337: ff_rdata <= 8'hB8;
			14'd1338: ff_rdata <= 8'h88;
			14'd1339: ff_rdata <= 8'h88;
			14'd1340: ff_rdata <= 8'h70;
			14'd1341: ff_rdata <= 8'h00;
			14'd1342: ff_rdata <= 8'h88;
			14'd1343: ff_rdata <= 8'h88;
			14'd1344: ff_rdata <= 8'h88;
			14'd1345: ff_rdata <= 8'hF8;
			14'd1346: ff_rdata <= 8'h88;
			14'd1347: ff_rdata <= 8'h88;
			14'd1348: ff_rdata <= 8'h88;
			14'd1349: ff_rdata <= 8'h00;
			14'd1350: ff_rdata <= 8'h70;
			14'd1351: ff_rdata <= 8'h20;
			14'd1352: ff_rdata <= 8'h20;
			14'd1353: ff_rdata <= 8'h20;
			14'd1354: ff_rdata <= 8'h20;
			14'd1355: ff_rdata <= 8'h20;
			14'd1356: ff_rdata <= 8'h70;
			14'd1357: ff_rdata <= 8'h00;
			14'd1358: ff_rdata <= 8'h38;
			14'd1359: ff_rdata <= 8'h10;
			14'd1360: ff_rdata <= 8'h10;
			14'd1361: ff_rdata <= 8'h10;
			14'd1362: ff_rdata <= 8'h90;
			14'd1363: ff_rdata <= 8'h90;
			14'd1364: ff_rdata <= 8'h60;
			14'd1365: ff_rdata <= 8'h00;
			14'd1366: ff_rdata <= 8'h88;
			14'd1367: ff_rdata <= 8'h90;
			14'd1368: ff_rdata <= 8'hA0;
			14'd1369: ff_rdata <= 8'hC0;
			14'd1370: ff_rdata <= 8'hA0;
			14'd1371: ff_rdata <= 8'h90;
			14'd1372: ff_rdata <= 8'h88;
			14'd1373: ff_rdata <= 8'h00;
			14'd1374: ff_rdata <= 8'h80;
			14'd1375: ff_rdata <= 8'h80;
			14'd1376: ff_rdata <= 8'h80;
			14'd1377: ff_rdata <= 8'h80;
			14'd1378: ff_rdata <= 8'h80;
			14'd1379: ff_rdata <= 8'h80;
			14'd1380: ff_rdata <= 8'hF8;
			14'd1381: ff_rdata <= 8'h00;
			14'd1382: ff_rdata <= 8'h88;
			14'd1383: ff_rdata <= 8'hD8;
			14'd1384: ff_rdata <= 8'hA8;
			14'd1385: ff_rdata <= 8'hA8;
			14'd1386: ff_rdata <= 8'h88;
			14'd1387: ff_rdata <= 8'h88;
			14'd1388: ff_rdata <= 8'h88;
			14'd1389: ff_rdata <= 8'h00;
			14'd1390: ff_rdata <= 8'h88;
			14'd1391: ff_rdata <= 8'hC8;
			14'd1392: ff_rdata <= 8'hC8;
			14'd1393: ff_rdata <= 8'hA8;
			14'd1394: ff_rdata <= 8'h98;
			14'd1395: ff_rdata <= 8'h98;
			14'd1396: ff_rdata <= 8'h88;
			14'd1397: ff_rdata <= 8'h00;
			14'd1398: ff_rdata <= 8'h70;
			14'd1399: ff_rdata <= 8'h88;
			14'd1400: ff_rdata <= 8'h88;
			14'd1401: ff_rdata <= 8'h88;
			14'd1402: ff_rdata <= 8'h88;
			14'd1403: ff_rdata <= 8'h88;
			14'd1404: ff_rdata <= 8'h70;
			14'd1405: ff_rdata <= 8'h00;
			14'd1406: ff_rdata <= 8'hF0;
			14'd1407: ff_rdata <= 8'h88;
			14'd1408: ff_rdata <= 8'h88;
			14'd1409: ff_rdata <= 8'hF0;
			14'd1410: ff_rdata <= 8'h80;
			14'd1411: ff_rdata <= 8'h80;
			14'd1412: ff_rdata <= 8'h80;
			14'd1413: ff_rdata <= 8'h00;
			14'd1414: ff_rdata <= 8'h70;
			14'd1415: ff_rdata <= 8'h88;
			14'd1416: ff_rdata <= 8'h88;
			14'd1417: ff_rdata <= 8'h88;
			14'd1418: ff_rdata <= 8'hA8;
			14'd1419: ff_rdata <= 8'h90;
			14'd1420: ff_rdata <= 8'h68;
			14'd1421: ff_rdata <= 8'h00;
			14'd1422: ff_rdata <= 8'hF0;
			14'd1423: ff_rdata <= 8'h88;
			14'd1424: ff_rdata <= 8'h88;
			14'd1425: ff_rdata <= 8'hF0;
			14'd1426: ff_rdata <= 8'hA0;
			14'd1427: ff_rdata <= 8'h90;
			14'd1428: ff_rdata <= 8'h88;
			14'd1429: ff_rdata <= 8'h00;
			14'd1430: ff_rdata <= 8'h70;
			14'd1431: ff_rdata <= 8'h88;
			14'd1432: ff_rdata <= 8'h80;
			14'd1433: ff_rdata <= 8'h70;
			14'd1434: ff_rdata <= 8'h08;
			14'd1435: ff_rdata <= 8'h88;
			14'd1436: ff_rdata <= 8'h70;
			14'd1437: ff_rdata <= 8'h00;
			14'd1438: ff_rdata <= 8'hF8;
			14'd1439: ff_rdata <= 8'h20;
			14'd1440: ff_rdata <= 8'h20;
			14'd1441: ff_rdata <= 8'h20;
			14'd1442: ff_rdata <= 8'h20;
			14'd1443: ff_rdata <= 8'h20;
			14'd1444: ff_rdata <= 8'h20;
			14'd1445: ff_rdata <= 8'h00;
			14'd1446: ff_rdata <= 8'h88;
			14'd1447: ff_rdata <= 8'h88;
			14'd1448: ff_rdata <= 8'h88;
			14'd1449: ff_rdata <= 8'h88;
			14'd1450: ff_rdata <= 8'h88;
			14'd1451: ff_rdata <= 8'h88;
			14'd1452: ff_rdata <= 8'h70;
			14'd1453: ff_rdata <= 8'h00;
			14'd1454: ff_rdata <= 8'h88;
			14'd1455: ff_rdata <= 8'h88;
			14'd1456: ff_rdata <= 8'h88;
			14'd1457: ff_rdata <= 8'h88;
			14'd1458: ff_rdata <= 8'h50;
			14'd1459: ff_rdata <= 8'h50;
			14'd1460: ff_rdata <= 8'h20;
			14'd1461: ff_rdata <= 8'h00;
			14'd1462: ff_rdata <= 8'h88;
			14'd1463: ff_rdata <= 8'h88;
			14'd1464: ff_rdata <= 8'h88;
			14'd1465: ff_rdata <= 8'hA8;
			14'd1466: ff_rdata <= 8'hA8;
			14'd1467: ff_rdata <= 8'hD8;
			14'd1468: ff_rdata <= 8'h88;
			14'd1469: ff_rdata <= 8'h00;
			14'd1470: ff_rdata <= 8'h88;
			14'd1471: ff_rdata <= 8'h88;
			14'd1472: ff_rdata <= 8'h50;
			14'd1473: ff_rdata <= 8'h20;
			14'd1474: ff_rdata <= 8'h50;
			14'd1475: ff_rdata <= 8'h88;
			14'd1476: ff_rdata <= 8'h88;
			14'd1477: ff_rdata <= 8'h00;
			14'd1478: ff_rdata <= 8'h88;
			14'd1479: ff_rdata <= 8'h88;
			14'd1480: ff_rdata <= 8'h88;
			14'd1481: ff_rdata <= 8'h70;
			14'd1482: ff_rdata <= 8'h20;
			14'd1483: ff_rdata <= 8'h20;
			14'd1484: ff_rdata <= 8'h20;
			14'd1485: ff_rdata <= 8'h00;
			14'd1486: ff_rdata <= 8'hF8;
			14'd1487: ff_rdata <= 8'h08;
			14'd1488: ff_rdata <= 8'h10;
			14'd1489: ff_rdata <= 8'h20;
			14'd1490: ff_rdata <= 8'h40;
			14'd1491: ff_rdata <= 8'h80;
			14'd1492: ff_rdata <= 8'hF8;
			14'd1493: ff_rdata <= 8'h00;
			14'd1494: ff_rdata <= 8'h70;
			14'd1495: ff_rdata <= 8'h40;
			14'd1496: ff_rdata <= 8'h40;
			14'd1497: ff_rdata <= 8'h40;
			14'd1498: ff_rdata <= 8'h40;
			14'd1499: ff_rdata <= 8'h40;
			14'd1500: ff_rdata <= 8'h70;
			14'd1501: ff_rdata <= 8'h00;
			14'd1502: ff_rdata <= 8'h88;
			14'd1503: ff_rdata <= 8'h50;
			14'd1504: ff_rdata <= 8'h20;
			14'd1505: ff_rdata <= 8'h70;
			14'd1506: ff_rdata <= 8'h20;
			14'd1507: ff_rdata <= 8'h70;
			14'd1508: ff_rdata <= 8'h20;
			14'd1509: ff_rdata <= 8'h00;
			14'd1510: ff_rdata <= 8'h70;
			14'd1511: ff_rdata <= 8'h10;
			14'd1512: ff_rdata <= 8'h10;
			14'd1513: ff_rdata <= 8'h10;
			14'd1514: ff_rdata <= 8'h10;
			14'd1515: ff_rdata <= 8'h10;
			14'd1516: ff_rdata <= 8'h70;
			14'd1517: ff_rdata <= 8'h00;
			14'd1518: ff_rdata <= 8'h20;
			14'd1519: ff_rdata <= 8'h50;
			14'd1520: ff_rdata <= 8'h88;
			14'd1521: ff_rdata <= 8'h00;
			14'd1522: ff_rdata <= 8'h00;
			14'd1523: ff_rdata <= 8'h00;
			14'd1524: ff_rdata <= 8'h00;
			14'd1525: ff_rdata <= 8'h00;
			14'd1526: ff_rdata <= 8'h00;
			14'd1527: ff_rdata <= 8'h00;
			14'd1528: ff_rdata <= 8'h00;
			14'd1529: ff_rdata <= 8'h00;
			14'd1530: ff_rdata <= 8'h00;
			14'd1531: ff_rdata <= 8'h00;
			14'd1532: ff_rdata <= 8'hF8;
			14'd1533: ff_rdata <= 8'h00;
			14'd1534: ff_rdata <= 8'h40;
			14'd1535: ff_rdata <= 8'h20;
			14'd1536: ff_rdata <= 8'h10;
			14'd1537: ff_rdata <= 8'h00;
			14'd1538: ff_rdata <= 8'h00;
			14'd1539: ff_rdata <= 8'h00;
			14'd1540: ff_rdata <= 8'h00;
			14'd1541: ff_rdata <= 8'h00;
			14'd1542: ff_rdata <= 8'h00;
			14'd1543: ff_rdata <= 8'h00;
			14'd1544: ff_rdata <= 8'h70;
			14'd1545: ff_rdata <= 8'h08;
			14'd1546: ff_rdata <= 8'h78;
			14'd1547: ff_rdata <= 8'h88;
			14'd1548: ff_rdata <= 8'h78;
			14'd1549: ff_rdata <= 8'h00;
			14'd1550: ff_rdata <= 8'h80;
			14'd1551: ff_rdata <= 8'h80;
			14'd1552: ff_rdata <= 8'hB0;
			14'd1553: ff_rdata <= 8'hC8;
			14'd1554: ff_rdata <= 8'h88;
			14'd1555: ff_rdata <= 8'hC8;
			14'd1556: ff_rdata <= 8'hB0;
			14'd1557: ff_rdata <= 8'h00;
			14'd1558: ff_rdata <= 8'h00;
			14'd1559: ff_rdata <= 8'h00;
			14'd1560: ff_rdata <= 8'h70;
			14'd1561: ff_rdata <= 8'h88;
			14'd1562: ff_rdata <= 8'h80;
			14'd1563: ff_rdata <= 8'h88;
			14'd1564: ff_rdata <= 8'h70;
			14'd1565: ff_rdata <= 8'h00;
			14'd1566: ff_rdata <= 8'h08;
			14'd1567: ff_rdata <= 8'h08;
			14'd1568: ff_rdata <= 8'h68;
			14'd1569: ff_rdata <= 8'h98;
			14'd1570: ff_rdata <= 8'h88;
			14'd1571: ff_rdata <= 8'h98;
			14'd1572: ff_rdata <= 8'h68;
			14'd1573: ff_rdata <= 8'h00;
			14'd1574: ff_rdata <= 8'h00;
			14'd1575: ff_rdata <= 8'h00;
			14'd1576: ff_rdata <= 8'h70;
			14'd1577: ff_rdata <= 8'h88;
			14'd1578: ff_rdata <= 8'hF8;
			14'd1579: ff_rdata <= 8'h80;
			14'd1580: ff_rdata <= 8'h70;
			14'd1581: ff_rdata <= 8'h00;
			14'd1582: ff_rdata <= 8'h10;
			14'd1583: ff_rdata <= 8'h28;
			14'd1584: ff_rdata <= 8'h20;
			14'd1585: ff_rdata <= 8'hF8;
			14'd1586: ff_rdata <= 8'h20;
			14'd1587: ff_rdata <= 8'h20;
			14'd1588: ff_rdata <= 8'h20;
			14'd1589: ff_rdata <= 8'h00;
			14'd1590: ff_rdata <= 8'h00;
			14'd1591: ff_rdata <= 8'h00;
			14'd1592: ff_rdata <= 8'h68;
			14'd1593: ff_rdata <= 8'h98;
			14'd1594: ff_rdata <= 8'h98;
			14'd1595: ff_rdata <= 8'h68;
			14'd1596: ff_rdata <= 8'h08;
			14'd1597: ff_rdata <= 8'h70;
			14'd1598: ff_rdata <= 8'h80;
			14'd1599: ff_rdata <= 8'h80;
			14'd1600: ff_rdata <= 8'hF0;
			14'd1601: ff_rdata <= 8'h88;
			14'd1602: ff_rdata <= 8'h88;
			14'd1603: ff_rdata <= 8'h88;
			14'd1604: ff_rdata <= 8'h88;
			14'd1605: ff_rdata <= 8'h00;
			14'd1606: ff_rdata <= 8'h20;
			14'd1607: ff_rdata <= 8'h00;
			14'd1608: ff_rdata <= 8'h60;
			14'd1609: ff_rdata <= 8'h20;
			14'd1610: ff_rdata <= 8'h20;
			14'd1611: ff_rdata <= 8'h20;
			14'd1612: ff_rdata <= 8'h70;
			14'd1613: ff_rdata <= 8'h00;
			14'd1614: ff_rdata <= 8'h10;
			14'd1615: ff_rdata <= 8'h00;
			14'd1616: ff_rdata <= 8'h30;
			14'd1617: ff_rdata <= 8'h10;
			14'd1618: ff_rdata <= 8'h10;
			14'd1619: ff_rdata <= 8'h10;
			14'd1620: ff_rdata <= 8'h90;
			14'd1621: ff_rdata <= 8'h60;
			14'd1622: ff_rdata <= 8'h40;
			14'd1623: ff_rdata <= 8'h40;
			14'd1624: ff_rdata <= 8'h48;
			14'd1625: ff_rdata <= 8'h50;
			14'd1626: ff_rdata <= 8'h60;
			14'd1627: ff_rdata <= 8'h50;
			14'd1628: ff_rdata <= 8'h48;
			14'd1629: ff_rdata <= 8'h00;
			14'd1630: ff_rdata <= 8'h60;
			14'd1631: ff_rdata <= 8'h20;
			14'd1632: ff_rdata <= 8'h20;
			14'd1633: ff_rdata <= 8'h20;
			14'd1634: ff_rdata <= 8'h20;
			14'd1635: ff_rdata <= 8'h20;
			14'd1636: ff_rdata <= 8'h70;
			14'd1637: ff_rdata <= 8'h00;
			14'd1638: ff_rdata <= 8'h00;
			14'd1639: ff_rdata <= 8'h00;
			14'd1640: ff_rdata <= 8'hD0;
			14'd1641: ff_rdata <= 8'hA8;
			14'd1642: ff_rdata <= 8'hA8;
			14'd1643: ff_rdata <= 8'hA8;
			14'd1644: ff_rdata <= 8'hA8;
			14'd1645: ff_rdata <= 8'h00;
			14'd1646: ff_rdata <= 8'h00;
			14'd1647: ff_rdata <= 8'h00;
			14'd1648: ff_rdata <= 8'hB0;
			14'd1649: ff_rdata <= 8'hC8;
			14'd1650: ff_rdata <= 8'h88;
			14'd1651: ff_rdata <= 8'h88;
			14'd1652: ff_rdata <= 8'h88;
			14'd1653: ff_rdata <= 8'h00;
			14'd1654: ff_rdata <= 8'h00;
			14'd1655: ff_rdata <= 8'h00;
			14'd1656: ff_rdata <= 8'h70;
			14'd1657: ff_rdata <= 8'h88;
			14'd1658: ff_rdata <= 8'h88;
			14'd1659: ff_rdata <= 8'h88;
			14'd1660: ff_rdata <= 8'h70;
			14'd1661: ff_rdata <= 8'h00;
			14'd1662: ff_rdata <= 8'h00;
			14'd1663: ff_rdata <= 8'h00;
			14'd1664: ff_rdata <= 8'hB0;
			14'd1665: ff_rdata <= 8'hC8;
			14'd1666: ff_rdata <= 8'hC8;
			14'd1667: ff_rdata <= 8'hB0;
			14'd1668: ff_rdata <= 8'h80;
			14'd1669: ff_rdata <= 8'h80;
			14'd1670: ff_rdata <= 8'h00;
			14'd1671: ff_rdata <= 8'h00;
			14'd1672: ff_rdata <= 8'h68;
			14'd1673: ff_rdata <= 8'h98;
			14'd1674: ff_rdata <= 8'h98;
			14'd1675: ff_rdata <= 8'h68;
			14'd1676: ff_rdata <= 8'h08;
			14'd1677: ff_rdata <= 8'h08;
			14'd1678: ff_rdata <= 8'h00;
			14'd1679: ff_rdata <= 8'h00;
			14'd1680: ff_rdata <= 8'hB0;
			14'd1681: ff_rdata <= 8'hC8;
			14'd1682: ff_rdata <= 8'h80;
			14'd1683: ff_rdata <= 8'h80;
			14'd1684: ff_rdata <= 8'h80;
			14'd1685: ff_rdata <= 8'h00;
			14'd1686: ff_rdata <= 8'h00;
			14'd1687: ff_rdata <= 8'h00;
			14'd1688: ff_rdata <= 8'h78;
			14'd1689: ff_rdata <= 8'h80;
			14'd1690: ff_rdata <= 8'hF0;
			14'd1691: ff_rdata <= 8'h08;
			14'd1692: ff_rdata <= 8'hF0;
			14'd1693: ff_rdata <= 8'h00;
			14'd1694: ff_rdata <= 8'h40;
			14'd1695: ff_rdata <= 8'h40;
			14'd1696: ff_rdata <= 8'hF0;
			14'd1697: ff_rdata <= 8'h40;
			14'd1698: ff_rdata <= 8'h40;
			14'd1699: ff_rdata <= 8'h48;
			14'd1700: ff_rdata <= 8'h30;
			14'd1701: ff_rdata <= 8'h00;
			14'd1702: ff_rdata <= 8'h00;
			14'd1703: ff_rdata <= 8'h00;
			14'd1704: ff_rdata <= 8'h90;
			14'd1705: ff_rdata <= 8'h90;
			14'd1706: ff_rdata <= 8'h90;
			14'd1707: ff_rdata <= 8'h90;
			14'd1708: ff_rdata <= 8'h68;
			14'd1709: ff_rdata <= 8'h00;
			14'd1710: ff_rdata <= 8'h00;
			14'd1711: ff_rdata <= 8'h00;
			14'd1712: ff_rdata <= 8'h88;
			14'd1713: ff_rdata <= 8'h88;
			14'd1714: ff_rdata <= 8'h88;
			14'd1715: ff_rdata <= 8'h50;
			14'd1716: ff_rdata <= 8'h20;
			14'd1717: ff_rdata <= 8'h00;
			14'd1718: ff_rdata <= 8'h00;
			14'd1719: ff_rdata <= 8'h00;
			14'd1720: ff_rdata <= 8'h88;
			14'd1721: ff_rdata <= 8'hA8;
			14'd1722: ff_rdata <= 8'hA8;
			14'd1723: ff_rdata <= 8'hA8;
			14'd1724: ff_rdata <= 8'h50;
			14'd1725: ff_rdata <= 8'h00;
			14'd1726: ff_rdata <= 8'h00;
			14'd1727: ff_rdata <= 8'h00;
			14'd1728: ff_rdata <= 8'h88;
			14'd1729: ff_rdata <= 8'h50;
			14'd1730: ff_rdata <= 8'h20;
			14'd1731: ff_rdata <= 8'h50;
			14'd1732: ff_rdata <= 8'h88;
			14'd1733: ff_rdata <= 8'h00;
			14'd1734: ff_rdata <= 8'h00;
			14'd1735: ff_rdata <= 8'h00;
			14'd1736: ff_rdata <= 8'h88;
			14'd1737: ff_rdata <= 8'h88;
			14'd1738: ff_rdata <= 8'h98;
			14'd1739: ff_rdata <= 8'h68;
			14'd1740: ff_rdata <= 8'h08;
			14'd1741: ff_rdata <= 8'h70;
			14'd1742: ff_rdata <= 8'h00;
			14'd1743: ff_rdata <= 8'h00;
			14'd1744: ff_rdata <= 8'hF8;
			14'd1745: ff_rdata <= 8'h10;
			14'd1746: ff_rdata <= 8'h20;
			14'd1747: ff_rdata <= 8'h40;
			14'd1748: ff_rdata <= 8'hF8;
			14'd1749: ff_rdata <= 8'h00;
			14'd1750: ff_rdata <= 8'h18;
			14'd1751: ff_rdata <= 8'h20;
			14'd1752: ff_rdata <= 8'h20;
			14'd1753: ff_rdata <= 8'h40;
			14'd1754: ff_rdata <= 8'h20;
			14'd1755: ff_rdata <= 8'h20;
			14'd1756: ff_rdata <= 8'h18;
			14'd1757: ff_rdata <= 8'h00;
			14'd1758: ff_rdata <= 8'h20;
			14'd1759: ff_rdata <= 8'h20;
			14'd1760: ff_rdata <= 8'h20;
			14'd1761: ff_rdata <= 8'h00;
			14'd1762: ff_rdata <= 8'h20;
			14'd1763: ff_rdata <= 8'h20;
			14'd1764: ff_rdata <= 8'h20;
			14'd1765: ff_rdata <= 8'h00;
			14'd1766: ff_rdata <= 8'hC0;
			14'd1767: ff_rdata <= 8'h20;
			14'd1768: ff_rdata <= 8'h20;
			14'd1769: ff_rdata <= 8'h10;
			14'd1770: ff_rdata <= 8'h20;
			14'd1771: ff_rdata <= 8'h20;
			14'd1772: ff_rdata <= 8'hC0;
			14'd1773: ff_rdata <= 8'h00;
			14'd1774: ff_rdata <= 8'h40;
			14'd1775: ff_rdata <= 8'hA8;
			14'd1776: ff_rdata <= 8'h10;
			14'd1777: ff_rdata <= 8'h00;
			14'd1778: ff_rdata <= 8'h00;
			14'd1779: ff_rdata <= 8'h00;
			14'd1780: ff_rdata <= 8'h00;
			14'd1781: ff_rdata <= 8'h00;
			14'd1782: ff_rdata <= 8'h00;
			14'd1783: ff_rdata <= 8'h00;
			14'd1784: ff_rdata <= 8'h00;
			14'd1785: ff_rdata <= 8'h00;
			14'd1786: ff_rdata <= 8'h00;
			14'd1787: ff_rdata <= 8'h00;
			14'd1788: ff_rdata <= 8'h00;
			14'd1789: ff_rdata <= 8'h00;
			14'd1790: ff_rdata <= 8'h10;
			14'd1791: ff_rdata <= 8'h38;
			14'd1792: ff_rdata <= 8'h7C;
			14'd1793: ff_rdata <= 8'hFE;
			14'd1794: ff_rdata <= 8'hFE;
			14'd1795: ff_rdata <= 8'h38;
			14'd1796: ff_rdata <= 8'h7C;
			14'd1797: ff_rdata <= 8'h00;
			14'd1798: ff_rdata <= 8'h6C;
			14'd1799: ff_rdata <= 8'hFE;
			14'd1800: ff_rdata <= 8'hFE;
			14'd1801: ff_rdata <= 8'hFE;
			14'd1802: ff_rdata <= 8'h7C;
			14'd1803: ff_rdata <= 8'h38;
			14'd1804: ff_rdata <= 8'h10;
			14'd1805: ff_rdata <= 8'h00;
			14'd1806: ff_rdata <= 8'h38;
			14'd1807: ff_rdata <= 8'h38;
			14'd1808: ff_rdata <= 8'hFE;
			14'd1809: ff_rdata <= 8'hFE;
			14'd1810: ff_rdata <= 8'hD6;
			14'd1811: ff_rdata <= 8'h10;
			14'd1812: ff_rdata <= 8'h7C;
			14'd1813: ff_rdata <= 8'h00;
			14'd1814: ff_rdata <= 8'h10;
			14'd1815: ff_rdata <= 8'h38;
			14'd1816: ff_rdata <= 8'h7C;
			14'd1817: ff_rdata <= 8'hFE;
			14'd1818: ff_rdata <= 8'h7C;
			14'd1819: ff_rdata <= 8'h38;
			14'd1820: ff_rdata <= 8'h10;
			14'd1821: ff_rdata <= 8'h00;
			14'd1822: ff_rdata <= 8'h00;
			14'd1823: ff_rdata <= 8'h78;
			14'd1824: ff_rdata <= 8'h84;
			14'd1825: ff_rdata <= 8'h84;
			14'd1826: ff_rdata <= 8'h84;
			14'd1827: ff_rdata <= 8'h84;
			14'd1828: ff_rdata <= 8'h78;
			14'd1829: ff_rdata <= 8'h00;
			14'd1830: ff_rdata <= 8'h00;
			14'd1831: ff_rdata <= 8'h78;
			14'd1832: ff_rdata <= 8'hFC;
			14'd1833: ff_rdata <= 8'hFC;
			14'd1834: ff_rdata <= 8'hFC;
			14'd1835: ff_rdata <= 8'hFC;
			14'd1836: ff_rdata <= 8'h78;
			14'd1837: ff_rdata <= 8'h00;
			14'd1838: ff_rdata <= 8'h20;
			14'd1839: ff_rdata <= 8'hF0;
			14'd1840: ff_rdata <= 8'h4C;
			14'd1841: ff_rdata <= 8'h70;
			14'd1842: ff_rdata <= 8'hA8;
			14'd1843: ff_rdata <= 8'h40;
			14'd1844: ff_rdata <= 8'h3C;
			14'd1845: ff_rdata <= 8'h00;
			14'd1846: ff_rdata <= 8'h00;
			14'd1847: ff_rdata <= 8'h20;
			14'd1848: ff_rdata <= 8'h78;
			14'd1849: ff_rdata <= 8'h20;
			14'd1850: ff_rdata <= 8'h78;
			14'd1851: ff_rdata <= 8'hB4;
			14'd1852: ff_rdata <= 8'h64;
			14'd1853: ff_rdata <= 8'h00;
			14'd1854: ff_rdata <= 8'h00;
			14'd1855: ff_rdata <= 8'h00;
			14'd1856: ff_rdata <= 8'h88;
			14'd1857: ff_rdata <= 8'h84;
			14'd1858: ff_rdata <= 8'h84;
			14'd1859: ff_rdata <= 8'h84;
			14'd1860: ff_rdata <= 8'h40;
			14'd1861: ff_rdata <= 8'h00;
			14'd1862: ff_rdata <= 8'h00;
			14'd1863: ff_rdata <= 8'h70;
			14'd1864: ff_rdata <= 8'h00;
			14'd1865: ff_rdata <= 8'h70;
			14'd1866: ff_rdata <= 8'h88;
			14'd1867: ff_rdata <= 8'h08;
			14'd1868: ff_rdata <= 8'h30;
			14'd1869: ff_rdata <= 8'h00;
			14'd1870: ff_rdata <= 8'h00;
			14'd1871: ff_rdata <= 8'h70;
			14'd1872: ff_rdata <= 8'h00;
			14'd1873: ff_rdata <= 8'hF0;
			14'd1874: ff_rdata <= 8'h20;
			14'd1875: ff_rdata <= 8'h60;
			14'd1876: ff_rdata <= 8'h98;
			14'd1877: ff_rdata <= 8'h00;
			14'd1878: ff_rdata <= 8'h00;
			14'd1879: ff_rdata <= 8'h20;
			14'd1880: ff_rdata <= 8'hF8;
			14'd1881: ff_rdata <= 8'h24;
			14'd1882: ff_rdata <= 8'h78;
			14'd1883: ff_rdata <= 8'hA4;
			14'd1884: ff_rdata <= 8'h68;
			14'd1885: ff_rdata <= 8'h00;
			14'd1886: ff_rdata <= 8'h00;
			14'd1887: ff_rdata <= 8'h90;
			14'd1888: ff_rdata <= 8'h58;
			14'd1889: ff_rdata <= 8'h64;
			14'd1890: ff_rdata <= 8'hA8;
			14'd1891: ff_rdata <= 8'h20;
			14'd1892: ff_rdata <= 8'h10;
			14'd1893: ff_rdata <= 8'h00;
			14'd1894: ff_rdata <= 8'h00;
			14'd1895: ff_rdata <= 8'h10;
			14'd1896: ff_rdata <= 8'hB8;
			14'd1897: ff_rdata <= 8'hD4;
			14'd1898: ff_rdata <= 8'h94;
			14'd1899: ff_rdata <= 8'h18;
			14'd1900: ff_rdata <= 8'h20;
			14'd1901: ff_rdata <= 8'h00;
			14'd1902: ff_rdata <= 8'h00;
			14'd1903: ff_rdata <= 8'h10;
			14'd1904: ff_rdata <= 8'h1C;
			14'd1905: ff_rdata <= 8'h10;
			14'd1906: ff_rdata <= 8'h70;
			14'd1907: ff_rdata <= 8'h98;
			14'd1908: ff_rdata <= 8'h74;
			14'd1909: ff_rdata <= 8'h00;
			14'd1910: ff_rdata <= 8'h00;
			14'd1911: ff_rdata <= 8'h00;
			14'd1912: ff_rdata <= 8'h00;
			14'd1913: ff_rdata <= 8'h78;
			14'd1914: ff_rdata <= 8'h04;
			14'd1915: ff_rdata <= 8'h04;
			14'd1916: ff_rdata <= 8'h38;
			14'd1917: ff_rdata <= 8'h00;
			14'd1918: ff_rdata <= 8'h00;
			14'd1919: ff_rdata <= 8'h00;
			14'd1920: ff_rdata <= 8'h00;
			14'd1921: ff_rdata <= 8'h00;
			14'd1922: ff_rdata <= 8'h00;
			14'd1923: ff_rdata <= 8'h00;
			14'd1924: ff_rdata <= 8'h00;
			14'd1925: ff_rdata <= 8'h00;
			14'd1926: ff_rdata <= 8'h20;
			14'd1927: ff_rdata <= 8'h7C;
			14'd1928: ff_rdata <= 8'h20;
			14'd1929: ff_rdata <= 8'h7C;
			14'd1930: ff_rdata <= 8'hAA;
			14'd1931: ff_rdata <= 8'h92;
			14'd1932: ff_rdata <= 8'h64;
			14'd1933: ff_rdata <= 8'h00;
			14'd1934: ff_rdata <= 8'h00;
			14'd1935: ff_rdata <= 8'h84;
			14'd1936: ff_rdata <= 8'h82;
			14'd1937: ff_rdata <= 8'h82;
			14'd1938: ff_rdata <= 8'h82;
			14'd1939: ff_rdata <= 8'h80;
			14'd1940: ff_rdata <= 8'h40;
			14'd1941: ff_rdata <= 8'h00;
			14'd1942: ff_rdata <= 8'h38;
			14'd1943: ff_rdata <= 8'h00;
			14'd1944: ff_rdata <= 8'h38;
			14'd1945: ff_rdata <= 8'h44;
			14'd1946: ff_rdata <= 8'h04;
			14'd1947: ff_rdata <= 8'h08;
			14'd1948: ff_rdata <= 8'h30;
			14'd1949: ff_rdata <= 8'h00;
			14'd1950: ff_rdata <= 8'h70;
			14'd1951: ff_rdata <= 8'h00;
			14'd1952: ff_rdata <= 8'hF8;
			14'd1953: ff_rdata <= 8'h10;
			14'd1954: ff_rdata <= 8'h20;
			14'd1955: ff_rdata <= 8'h60;
			14'd1956: ff_rdata <= 8'h9C;
			14'd1957: ff_rdata <= 8'h00;
			14'd1958: ff_rdata <= 8'h24;
			14'd1959: ff_rdata <= 8'hFA;
			14'd1960: ff_rdata <= 8'h20;
			14'd1961: ff_rdata <= 8'h7C;
			14'd1962: ff_rdata <= 8'hA2;
			14'd1963: ff_rdata <= 8'hA2;
			14'd1964: ff_rdata <= 8'h44;
			14'd1965: ff_rdata <= 8'h00;
			14'd1966: ff_rdata <= 8'h40;
			14'd1967: ff_rdata <= 8'h44;
			14'd1968: ff_rdata <= 8'hF2;
			14'd1969: ff_rdata <= 8'h4A;
			14'd1970: ff_rdata <= 8'h48;
			14'd1971: ff_rdata <= 8'h88;
			14'd1972: ff_rdata <= 8'h30;
			14'd1973: ff_rdata <= 8'h00;
			14'd1974: ff_rdata <= 8'h20;
			14'd1975: ff_rdata <= 8'hFC;
			14'd1976: ff_rdata <= 8'h10;
			14'd1977: ff_rdata <= 8'hFC;
			14'd1978: ff_rdata <= 8'h08;
			14'd1979: ff_rdata <= 8'h80;
			14'd1980: ff_rdata <= 8'h78;
			14'd1981: ff_rdata <= 8'h00;
			14'd1982: ff_rdata <= 8'h08;
			14'd1983: ff_rdata <= 8'h10;
			14'd1984: ff_rdata <= 8'h20;
			14'd1985: ff_rdata <= 8'h40;
			14'd1986: ff_rdata <= 8'h20;
			14'd1987: ff_rdata <= 8'h10;
			14'd1988: ff_rdata <= 8'h08;
			14'd1989: ff_rdata <= 8'h00;
			14'd1990: ff_rdata <= 8'h04;
			14'd1991: ff_rdata <= 8'h84;
			14'd1992: ff_rdata <= 8'h9E;
			14'd1993: ff_rdata <= 8'h84;
			14'd1994: ff_rdata <= 8'h84;
			14'd1995: ff_rdata <= 8'h84;
			14'd1996: ff_rdata <= 8'h48;
			14'd1997: ff_rdata <= 8'h00;
			14'd1998: ff_rdata <= 8'h78;
			14'd1999: ff_rdata <= 8'h04;
			14'd2000: ff_rdata <= 8'h00;
			14'd2001: ff_rdata <= 8'h00;
			14'd2002: ff_rdata <= 8'h00;
			14'd2003: ff_rdata <= 8'h80;
			14'd2004: ff_rdata <= 8'h7C;
			14'd2005: ff_rdata <= 8'h00;
			14'd2006: ff_rdata <= 8'h10;
			14'd2007: ff_rdata <= 8'hFE;
			14'd2008: ff_rdata <= 8'h08;
			14'd2009: ff_rdata <= 8'h04;
			14'd2010: ff_rdata <= 8'h04;
			14'd2011: ff_rdata <= 8'h80;
			14'd2012: ff_rdata <= 8'h78;
			14'd2013: ff_rdata <= 8'h00;
			14'd2014: ff_rdata <= 8'h80;
			14'd2015: ff_rdata <= 8'h80;
			14'd2016: ff_rdata <= 8'h80;
			14'd2017: ff_rdata <= 8'h80;
			14'd2018: ff_rdata <= 8'h84;
			14'd2019: ff_rdata <= 8'h88;
			14'd2020: ff_rdata <= 8'h70;
			14'd2021: ff_rdata <= 8'h00;
			14'd2022: ff_rdata <= 8'h08;
			14'd2023: ff_rdata <= 8'hFE;
			14'd2024: ff_rdata <= 8'h38;
			14'd2025: ff_rdata <= 8'h48;
			14'd2026: ff_rdata <= 8'h38;
			14'd2027: ff_rdata <= 8'h08;
			14'd2028: ff_rdata <= 8'h10;
			14'd2029: ff_rdata <= 8'h00;
			14'd2030: ff_rdata <= 8'h44;
			14'd2031: ff_rdata <= 8'h44;
			14'd2032: ff_rdata <= 8'hFE;
			14'd2033: ff_rdata <= 8'h44;
			14'd2034: ff_rdata <= 8'h48;
			14'd2035: ff_rdata <= 8'h40;
			14'd2036: ff_rdata <= 8'h3C;
			14'd2037: ff_rdata <= 8'h00;
			14'd2038: ff_rdata <= 8'h44;
			14'd2039: ff_rdata <= 8'h28;
			14'd2040: ff_rdata <= 8'hFE;
			14'd2041: ff_rdata <= 8'h20;
			14'd2042: ff_rdata <= 8'h40;
			14'd2043: ff_rdata <= 8'h40;
			14'd2044: ff_rdata <= 8'h3C;
			14'd2045: ff_rdata <= 8'h00;
			14'd2046: ff_rdata <= 8'h00;
			14'd2047: ff_rdata <= 8'h00;
			14'd2048: ff_rdata <= 8'h00;
			14'd2049: ff_rdata <= 8'h00;
			14'd2050: ff_rdata <= 8'h00;
			14'd2051: ff_rdata <= 8'h00;
			14'd2052: ff_rdata <= 8'h00;
			14'd2053: ff_rdata <= 8'h00;
			14'd2054: ff_rdata <= 8'h00;
			14'd2055: ff_rdata <= 8'h00;
			14'd2056: ff_rdata <= 8'h00;
			14'd2057: ff_rdata <= 8'h00;
			14'd2058: ff_rdata <= 8'h60;
			14'd2059: ff_rdata <= 8'h90;
			14'd2060: ff_rdata <= 8'h60;
			14'd2061: ff_rdata <= 8'h00;
			14'd2062: ff_rdata <= 8'h38;
			14'd2063: ff_rdata <= 8'h20;
			14'd2064: ff_rdata <= 8'h20;
			14'd2065: ff_rdata <= 8'h20;
			14'd2066: ff_rdata <= 8'h00;
			14'd2067: ff_rdata <= 8'h00;
			14'd2068: ff_rdata <= 8'h00;
			14'd2069: ff_rdata <= 8'h00;
			14'd2070: ff_rdata <= 8'h00;
			14'd2071: ff_rdata <= 8'h00;
			14'd2072: ff_rdata <= 8'h00;
			14'd2073: ff_rdata <= 8'h20;
			14'd2074: ff_rdata <= 8'h20;
			14'd2075: ff_rdata <= 8'h20;
			14'd2076: ff_rdata <= 8'hE0;
			14'd2077: ff_rdata <= 8'h00;
			14'd2078: ff_rdata <= 8'h00;
			14'd2079: ff_rdata <= 8'h00;
			14'd2080: ff_rdata <= 8'h00;
			14'd2081: ff_rdata <= 8'h00;
			14'd2082: ff_rdata <= 8'h80;
			14'd2083: ff_rdata <= 8'h40;
			14'd2084: ff_rdata <= 8'h20;
			14'd2085: ff_rdata <= 8'h00;
			14'd2086: ff_rdata <= 8'h00;
			14'd2087: ff_rdata <= 8'h00;
			14'd2088: ff_rdata <= 8'h00;
			14'd2089: ff_rdata <= 8'h30;
			14'd2090: ff_rdata <= 8'h30;
			14'd2091: ff_rdata <= 8'h00;
			14'd2092: ff_rdata <= 8'h00;
			14'd2093: ff_rdata <= 8'h00;
			14'd2094: ff_rdata <= 8'hF8;
			14'd2095: ff_rdata <= 8'h08;
			14'd2096: ff_rdata <= 8'hF8;
			14'd2097: ff_rdata <= 8'h08;
			14'd2098: ff_rdata <= 8'h10;
			14'd2099: ff_rdata <= 8'h20;
			14'd2100: ff_rdata <= 8'h40;
			14'd2101: ff_rdata <= 8'h00;
			14'd2102: ff_rdata <= 8'h00;
			14'd2103: ff_rdata <= 8'h00;
			14'd2104: ff_rdata <= 8'hF0;
			14'd2105: ff_rdata <= 8'h10;
			14'd2106: ff_rdata <= 8'h60;
			14'd2107: ff_rdata <= 8'h40;
			14'd2108: ff_rdata <= 8'h80;
			14'd2109: ff_rdata <= 8'h00;
			14'd2110: ff_rdata <= 8'h00;
			14'd2111: ff_rdata <= 8'h10;
			14'd2112: ff_rdata <= 8'h20;
			14'd2113: ff_rdata <= 8'h60;
			14'd2114: ff_rdata <= 8'hA0;
			14'd2115: ff_rdata <= 8'h20;
			14'd2116: ff_rdata <= 8'h20;
			14'd2117: ff_rdata <= 8'h00;
			14'd2118: ff_rdata <= 8'h00;
			14'd2119: ff_rdata <= 8'h20;
			14'd2120: ff_rdata <= 8'hF0;
			14'd2121: ff_rdata <= 8'h90;
			14'd2122: ff_rdata <= 8'h10;
			14'd2123: ff_rdata <= 8'h20;
			14'd2124: ff_rdata <= 8'h40;
			14'd2125: ff_rdata <= 8'h00;
			14'd2126: ff_rdata <= 8'h00;
			14'd2127: ff_rdata <= 8'h00;
			14'd2128: ff_rdata <= 8'hF0;
			14'd2129: ff_rdata <= 8'h20;
			14'd2130: ff_rdata <= 8'h20;
			14'd2131: ff_rdata <= 8'h20;
			14'd2132: ff_rdata <= 8'hF0;
			14'd2133: ff_rdata <= 8'h00;
			14'd2134: ff_rdata <= 8'h00;
			14'd2135: ff_rdata <= 8'h20;
			14'd2136: ff_rdata <= 8'hF0;
			14'd2137: ff_rdata <= 8'h60;
			14'd2138: ff_rdata <= 8'hA0;
			14'd2139: ff_rdata <= 8'hA0;
			14'd2140: ff_rdata <= 8'h20;
			14'd2141: ff_rdata <= 8'h00;
			14'd2142: ff_rdata <= 8'h00;
			14'd2143: ff_rdata <= 8'h40;
			14'd2144: ff_rdata <= 8'hF8;
			14'd2145: ff_rdata <= 8'h48;
			14'd2146: ff_rdata <= 8'h50;
			14'd2147: ff_rdata <= 8'h40;
			14'd2148: ff_rdata <= 8'h40;
			14'd2149: ff_rdata <= 8'h00;
			14'd2150: ff_rdata <= 8'h00;
			14'd2151: ff_rdata <= 8'h00;
			14'd2152: ff_rdata <= 8'h70;
			14'd2153: ff_rdata <= 8'h10;
			14'd2154: ff_rdata <= 8'h10;
			14'd2155: ff_rdata <= 8'h10;
			14'd2156: ff_rdata <= 8'hF8;
			14'd2157: ff_rdata <= 8'h00;
			14'd2158: ff_rdata <= 8'h00;
			14'd2159: ff_rdata <= 8'h00;
			14'd2160: ff_rdata <= 8'hF0;
			14'd2161: ff_rdata <= 8'h10;
			14'd2162: ff_rdata <= 8'hF0;
			14'd2163: ff_rdata <= 8'h10;
			14'd2164: ff_rdata <= 8'hF0;
			14'd2165: ff_rdata <= 8'h00;
			14'd2166: ff_rdata <= 8'h00;
			14'd2167: ff_rdata <= 8'h00;
			14'd2168: ff_rdata <= 8'hA8;
			14'd2169: ff_rdata <= 8'hA8;
			14'd2170: ff_rdata <= 8'h08;
			14'd2171: ff_rdata <= 8'h10;
			14'd2172: ff_rdata <= 8'h20;
			14'd2173: ff_rdata <= 8'h00;
			14'd2174: ff_rdata <= 8'h00;
			14'd2175: ff_rdata <= 8'h00;
			14'd2176: ff_rdata <= 8'h80;
			14'd2177: ff_rdata <= 8'h7C;
			14'd2178: ff_rdata <= 8'h00;
			14'd2179: ff_rdata <= 8'h00;
			14'd2180: ff_rdata <= 8'h00;
			14'd2181: ff_rdata <= 8'h00;
			14'd2182: ff_rdata <= 8'hF8;
			14'd2183: ff_rdata <= 8'h08;
			14'd2184: ff_rdata <= 8'h28;
			14'd2185: ff_rdata <= 8'h30;
			14'd2186: ff_rdata <= 8'h20;
			14'd2187: ff_rdata <= 8'h20;
			14'd2188: ff_rdata <= 8'h40;
			14'd2189: ff_rdata <= 8'h00;
			14'd2190: ff_rdata <= 8'h08;
			14'd2191: ff_rdata <= 8'h10;
			14'd2192: ff_rdata <= 8'h20;
			14'd2193: ff_rdata <= 8'h60;
			14'd2194: ff_rdata <= 8'hA0;
			14'd2195: ff_rdata <= 8'h20;
			14'd2196: ff_rdata <= 8'h20;
			14'd2197: ff_rdata <= 8'h00;
			14'd2198: ff_rdata <= 8'h20;
			14'd2199: ff_rdata <= 8'hF8;
			14'd2200: ff_rdata <= 8'h88;
			14'd2201: ff_rdata <= 8'h88;
			14'd2202: ff_rdata <= 8'h08;
			14'd2203: ff_rdata <= 8'h10;
			14'd2204: ff_rdata <= 8'h20;
			14'd2205: ff_rdata <= 8'h00;
			14'd2206: ff_rdata <= 8'h00;
			14'd2207: ff_rdata <= 8'hF8;
			14'd2208: ff_rdata <= 8'h20;
			14'd2209: ff_rdata <= 8'h20;
			14'd2210: ff_rdata <= 8'h20;
			14'd2211: ff_rdata <= 8'h20;
			14'd2212: ff_rdata <= 8'hF8;
			14'd2213: ff_rdata <= 8'h00;
			14'd2214: ff_rdata <= 8'h10;
			14'd2215: ff_rdata <= 8'hF8;
			14'd2216: ff_rdata <= 8'h10;
			14'd2217: ff_rdata <= 8'h30;
			14'd2218: ff_rdata <= 8'h50;
			14'd2219: ff_rdata <= 8'h90;
			14'd2220: ff_rdata <= 8'h10;
			14'd2221: ff_rdata <= 8'h00;
			14'd2222: ff_rdata <= 8'h20;
			14'd2223: ff_rdata <= 8'hF8;
			14'd2224: ff_rdata <= 8'h28;
			14'd2225: ff_rdata <= 8'h28;
			14'd2226: ff_rdata <= 8'h28;
			14'd2227: ff_rdata <= 8'h48;
			14'd2228: ff_rdata <= 8'h88;
			14'd2229: ff_rdata <= 8'h00;
			14'd2230: ff_rdata <= 8'h20;
			14'd2231: ff_rdata <= 8'hF8;
			14'd2232: ff_rdata <= 8'h20;
			14'd2233: ff_rdata <= 8'hF8;
			14'd2234: ff_rdata <= 8'h20;
			14'd2235: ff_rdata <= 8'h20;
			14'd2236: ff_rdata <= 8'h20;
			14'd2237: ff_rdata <= 8'h00;
			14'd2238: ff_rdata <= 8'h78;
			14'd2239: ff_rdata <= 8'h48;
			14'd2240: ff_rdata <= 8'h88;
			14'd2241: ff_rdata <= 8'h08;
			14'd2242: ff_rdata <= 8'h08;
			14'd2243: ff_rdata <= 8'h10;
			14'd2244: ff_rdata <= 8'h20;
			14'd2245: ff_rdata <= 8'h00;
			14'd2246: ff_rdata <= 8'h40;
			14'd2247: ff_rdata <= 8'h78;
			14'd2248: ff_rdata <= 8'h50;
			14'd2249: ff_rdata <= 8'h90;
			14'd2250: ff_rdata <= 8'h10;
			14'd2251: ff_rdata <= 8'h10;
			14'd2252: ff_rdata <= 8'h20;
			14'd2253: ff_rdata <= 8'h00;
			14'd2254: ff_rdata <= 8'h00;
			14'd2255: ff_rdata <= 8'hF8;
			14'd2256: ff_rdata <= 8'h08;
			14'd2257: ff_rdata <= 8'h08;
			14'd2258: ff_rdata <= 8'h08;
			14'd2259: ff_rdata <= 8'h08;
			14'd2260: ff_rdata <= 8'hF8;
			14'd2261: ff_rdata <= 8'h00;
			14'd2262: ff_rdata <= 8'h50;
			14'd2263: ff_rdata <= 8'hF8;
			14'd2264: ff_rdata <= 8'h50;
			14'd2265: ff_rdata <= 8'h50;
			14'd2266: ff_rdata <= 8'h10;
			14'd2267: ff_rdata <= 8'h10;
			14'd2268: ff_rdata <= 8'h20;
			14'd2269: ff_rdata <= 8'h00;
			14'd2270: ff_rdata <= 8'h00;
			14'd2271: ff_rdata <= 8'hC0;
			14'd2272: ff_rdata <= 8'h08;
			14'd2273: ff_rdata <= 8'hC8;
			14'd2274: ff_rdata <= 8'h08;
			14'd2275: ff_rdata <= 8'h10;
			14'd2276: ff_rdata <= 8'hE0;
			14'd2277: ff_rdata <= 8'h00;
			14'd2278: ff_rdata <= 8'h00;
			14'd2279: ff_rdata <= 8'hF8;
			14'd2280: ff_rdata <= 8'h08;
			14'd2281: ff_rdata <= 8'h10;
			14'd2282: ff_rdata <= 8'h20;
			14'd2283: ff_rdata <= 8'h50;
			14'd2284: ff_rdata <= 8'h88;
			14'd2285: ff_rdata <= 8'h00;
			14'd2286: ff_rdata <= 8'h40;
			14'd2287: ff_rdata <= 8'hF8;
			14'd2288: ff_rdata <= 8'h48;
			14'd2289: ff_rdata <= 8'h50;
			14'd2290: ff_rdata <= 8'h40;
			14'd2291: ff_rdata <= 8'h40;
			14'd2292: ff_rdata <= 8'h38;
			14'd2293: ff_rdata <= 8'h00;
			14'd2294: ff_rdata <= 8'h88;
			14'd2295: ff_rdata <= 8'h88;
			14'd2296: ff_rdata <= 8'h48;
			14'd2297: ff_rdata <= 8'h08;
			14'd2298: ff_rdata <= 8'h10;
			14'd2299: ff_rdata <= 8'h20;
			14'd2300: ff_rdata <= 8'h40;
			14'd2301: ff_rdata <= 8'h00;
			14'd2302: ff_rdata <= 8'h78;
			14'd2303: ff_rdata <= 8'h48;
			14'd2304: ff_rdata <= 8'h78;
			14'd2305: ff_rdata <= 8'h88;
			14'd2306: ff_rdata <= 8'h08;
			14'd2307: ff_rdata <= 8'h10;
			14'd2308: ff_rdata <= 8'h20;
			14'd2309: ff_rdata <= 8'h00;
			14'd2310: ff_rdata <= 8'h10;
			14'd2311: ff_rdata <= 8'hE0;
			14'd2312: ff_rdata <= 8'h20;
			14'd2313: ff_rdata <= 8'hF8;
			14'd2314: ff_rdata <= 8'h20;
			14'd2315: ff_rdata <= 8'h20;
			14'd2316: ff_rdata <= 8'h40;
			14'd2317: ff_rdata <= 8'h00;
			14'd2318: ff_rdata <= 8'hA8;
			14'd2319: ff_rdata <= 8'hA8;
			14'd2320: ff_rdata <= 8'hA8;
			14'd2321: ff_rdata <= 8'h08;
			14'd2322: ff_rdata <= 8'h08;
			14'd2323: ff_rdata <= 8'h10;
			14'd2324: ff_rdata <= 8'h20;
			14'd2325: ff_rdata <= 8'h00;
			14'd2326: ff_rdata <= 8'h70;
			14'd2327: ff_rdata <= 8'h00;
			14'd2328: ff_rdata <= 8'hF8;
			14'd2329: ff_rdata <= 8'h20;
			14'd2330: ff_rdata <= 8'h20;
			14'd2331: ff_rdata <= 8'h20;
			14'd2332: ff_rdata <= 8'h40;
			14'd2333: ff_rdata <= 8'h00;
			14'd2334: ff_rdata <= 8'h40;
			14'd2335: ff_rdata <= 8'h40;
			14'd2336: ff_rdata <= 8'h60;
			14'd2337: ff_rdata <= 8'h50;
			14'd2338: ff_rdata <= 8'h48;
			14'd2339: ff_rdata <= 8'h40;
			14'd2340: ff_rdata <= 8'h40;
			14'd2341: ff_rdata <= 8'h00;
			14'd2342: ff_rdata <= 8'h20;
			14'd2343: ff_rdata <= 8'hF8;
			14'd2344: ff_rdata <= 8'h20;
			14'd2345: ff_rdata <= 8'h20;
			14'd2346: ff_rdata <= 8'h20;
			14'd2347: ff_rdata <= 8'h20;
			14'd2348: ff_rdata <= 8'h40;
			14'd2349: ff_rdata <= 8'h00;
			14'd2350: ff_rdata <= 8'h00;
			14'd2351: ff_rdata <= 8'h70;
			14'd2352: ff_rdata <= 8'h00;
			14'd2353: ff_rdata <= 8'h00;
			14'd2354: ff_rdata <= 8'h00;
			14'd2355: ff_rdata <= 8'h00;
			14'd2356: ff_rdata <= 8'hF8;
			14'd2357: ff_rdata <= 8'h00;
			14'd2358: ff_rdata <= 8'h00;
			14'd2359: ff_rdata <= 8'hF8;
			14'd2360: ff_rdata <= 8'h08;
			14'd2361: ff_rdata <= 8'hD0;
			14'd2362: ff_rdata <= 8'h20;
			14'd2363: ff_rdata <= 8'h50;
			14'd2364: ff_rdata <= 8'h88;
			14'd2365: ff_rdata <= 8'h00;
			14'd2366: ff_rdata <= 8'h20;
			14'd2367: ff_rdata <= 8'hF8;
			14'd2368: ff_rdata <= 8'h08;
			14'd2369: ff_rdata <= 8'h30;
			14'd2370: ff_rdata <= 8'hE8;
			14'd2371: ff_rdata <= 8'h20;
			14'd2372: ff_rdata <= 8'h20;
			14'd2373: ff_rdata <= 8'h00;
			14'd2374: ff_rdata <= 8'h08;
			14'd2375: ff_rdata <= 8'h08;
			14'd2376: ff_rdata <= 8'h08;
			14'd2377: ff_rdata <= 8'h10;
			14'd2378: ff_rdata <= 8'h20;
			14'd2379: ff_rdata <= 8'h40;
			14'd2380: ff_rdata <= 8'h80;
			14'd2381: ff_rdata <= 8'h00;
			14'd2382: ff_rdata <= 8'h20;
			14'd2383: ff_rdata <= 8'h10;
			14'd2384: ff_rdata <= 8'h48;
			14'd2385: ff_rdata <= 8'h48;
			14'd2386: ff_rdata <= 8'h48;
			14'd2387: ff_rdata <= 8'h48;
			14'd2388: ff_rdata <= 8'h88;
			14'd2389: ff_rdata <= 8'h00;
			14'd2390: ff_rdata <= 8'h80;
			14'd2391: ff_rdata <= 8'h80;
			14'd2392: ff_rdata <= 8'hF8;
			14'd2393: ff_rdata <= 8'h80;
			14'd2394: ff_rdata <= 8'h80;
			14'd2395: ff_rdata <= 8'h80;
			14'd2396: ff_rdata <= 8'h78;
			14'd2397: ff_rdata <= 8'h00;
			14'd2398: ff_rdata <= 8'hF8;
			14'd2399: ff_rdata <= 8'h08;
			14'd2400: ff_rdata <= 8'h08;
			14'd2401: ff_rdata <= 8'h08;
			14'd2402: ff_rdata <= 8'h10;
			14'd2403: ff_rdata <= 8'h20;
			14'd2404: ff_rdata <= 8'h40;
			14'd2405: ff_rdata <= 8'h00;
			14'd2406: ff_rdata <= 8'h00;
			14'd2407: ff_rdata <= 8'h40;
			14'd2408: ff_rdata <= 8'hA0;
			14'd2409: ff_rdata <= 8'h10;
			14'd2410: ff_rdata <= 8'h08;
			14'd2411: ff_rdata <= 8'h08;
			14'd2412: ff_rdata <= 8'h00;
			14'd2413: ff_rdata <= 8'h00;
			14'd2414: ff_rdata <= 8'h20;
			14'd2415: ff_rdata <= 8'hF8;
			14'd2416: ff_rdata <= 8'h20;
			14'd2417: ff_rdata <= 8'h20;
			14'd2418: ff_rdata <= 8'hA8;
			14'd2419: ff_rdata <= 8'hA8;
			14'd2420: ff_rdata <= 8'h20;
			14'd2421: ff_rdata <= 8'h00;
			14'd2422: ff_rdata <= 8'h00;
			14'd2423: ff_rdata <= 8'hF8;
			14'd2424: ff_rdata <= 8'h08;
			14'd2425: ff_rdata <= 8'h08;
			14'd2426: ff_rdata <= 8'h50;
			14'd2427: ff_rdata <= 8'h20;
			14'd2428: ff_rdata <= 8'h10;
			14'd2429: ff_rdata <= 8'h00;
			14'd2430: ff_rdata <= 8'hF0;
			14'd2431: ff_rdata <= 8'h00;
			14'd2432: ff_rdata <= 8'h60;
			14'd2433: ff_rdata <= 8'h00;
			14'd2434: ff_rdata <= 8'h00;
			14'd2435: ff_rdata <= 8'hF0;
			14'd2436: ff_rdata <= 8'h08;
			14'd2437: ff_rdata <= 8'h00;
			14'd2438: ff_rdata <= 8'h10;
			14'd2439: ff_rdata <= 8'h20;
			14'd2440: ff_rdata <= 8'h40;
			14'd2441: ff_rdata <= 8'h80;
			14'd2442: ff_rdata <= 8'h90;
			14'd2443: ff_rdata <= 8'h88;
			14'd2444: ff_rdata <= 8'hF8;
			14'd2445: ff_rdata <= 8'h00;
			14'd2446: ff_rdata <= 8'h08;
			14'd2447: ff_rdata <= 8'h08;
			14'd2448: ff_rdata <= 8'h08;
			14'd2449: ff_rdata <= 8'h50;
			14'd2450: ff_rdata <= 8'h20;
			14'd2451: ff_rdata <= 8'h50;
			14'd2452: ff_rdata <= 8'h80;
			14'd2453: ff_rdata <= 8'h00;
			14'd2454: ff_rdata <= 8'h78;
			14'd2455: ff_rdata <= 8'h20;
			14'd2456: ff_rdata <= 8'hF8;
			14'd2457: ff_rdata <= 8'h20;
			14'd2458: ff_rdata <= 8'h20;
			14'd2459: ff_rdata <= 8'h20;
			14'd2460: ff_rdata <= 8'h18;
			14'd2461: ff_rdata <= 8'h00;
			14'd2462: ff_rdata <= 8'h40;
			14'd2463: ff_rdata <= 8'hF8;
			14'd2464: ff_rdata <= 8'h48;
			14'd2465: ff_rdata <= 8'h48;
			14'd2466: ff_rdata <= 8'h50;
			14'd2467: ff_rdata <= 8'h40;
			14'd2468: ff_rdata <= 8'h40;
			14'd2469: ff_rdata <= 8'h00;
			14'd2470: ff_rdata <= 8'h00;
			14'd2471: ff_rdata <= 8'h70;
			14'd2472: ff_rdata <= 8'h10;
			14'd2473: ff_rdata <= 8'h10;
			14'd2474: ff_rdata <= 8'h10;
			14'd2475: ff_rdata <= 8'h10;
			14'd2476: ff_rdata <= 8'hF8;
			14'd2477: ff_rdata <= 8'h00;
			14'd2478: ff_rdata <= 8'h00;
			14'd2479: ff_rdata <= 8'hF8;
			14'd2480: ff_rdata <= 8'h08;
			14'd2481: ff_rdata <= 8'hF8;
			14'd2482: ff_rdata <= 8'h08;
			14'd2483: ff_rdata <= 8'h08;
			14'd2484: ff_rdata <= 8'hF8;
			14'd2485: ff_rdata <= 8'h00;
			14'd2486: ff_rdata <= 8'h70;
			14'd2487: ff_rdata <= 8'h00;
			14'd2488: ff_rdata <= 8'hF8;
			14'd2489: ff_rdata <= 8'h08;
			14'd2490: ff_rdata <= 8'h08;
			14'd2491: ff_rdata <= 8'h10;
			14'd2492: ff_rdata <= 8'h20;
			14'd2493: ff_rdata <= 8'h00;
			14'd2494: ff_rdata <= 8'h48;
			14'd2495: ff_rdata <= 8'h48;
			14'd2496: ff_rdata <= 8'h48;
			14'd2497: ff_rdata <= 8'h48;
			14'd2498: ff_rdata <= 8'h48;
			14'd2499: ff_rdata <= 8'h10;
			14'd2500: ff_rdata <= 8'h20;
			14'd2501: ff_rdata <= 8'h00;
			14'd2502: ff_rdata <= 8'h10;
			14'd2503: ff_rdata <= 8'h50;
			14'd2504: ff_rdata <= 8'h50;
			14'd2505: ff_rdata <= 8'h50;
			14'd2506: ff_rdata <= 8'h50;
			14'd2507: ff_rdata <= 8'h58;
			14'd2508: ff_rdata <= 8'h90;
			14'd2509: ff_rdata <= 8'h00;
			14'd2510: ff_rdata <= 8'h40;
			14'd2511: ff_rdata <= 8'h40;
			14'd2512: ff_rdata <= 8'h40;
			14'd2513: ff_rdata <= 8'h48;
			14'd2514: ff_rdata <= 8'h48;
			14'd2515: ff_rdata <= 8'h50;
			14'd2516: ff_rdata <= 8'h60;
			14'd2517: ff_rdata <= 8'h00;
			14'd2518: ff_rdata <= 8'h00;
			14'd2519: ff_rdata <= 8'hF8;
			14'd2520: ff_rdata <= 8'h88;
			14'd2521: ff_rdata <= 8'h88;
			14'd2522: ff_rdata <= 8'h88;
			14'd2523: ff_rdata <= 8'h88;
			14'd2524: ff_rdata <= 8'hF8;
			14'd2525: ff_rdata <= 8'h00;
			14'd2526: ff_rdata <= 8'hF8;
			14'd2527: ff_rdata <= 8'h88;
			14'd2528: ff_rdata <= 8'h88;
			14'd2529: ff_rdata <= 8'h08;
			14'd2530: ff_rdata <= 8'h08;
			14'd2531: ff_rdata <= 8'h10;
			14'd2532: ff_rdata <= 8'h20;
			14'd2533: ff_rdata <= 8'h00;
			14'd2534: ff_rdata <= 8'h00;
			14'd2535: ff_rdata <= 8'hC0;
			14'd2536: ff_rdata <= 8'h00;
			14'd2537: ff_rdata <= 8'h08;
			14'd2538: ff_rdata <= 8'h08;
			14'd2539: ff_rdata <= 8'h10;
			14'd2540: ff_rdata <= 8'hE0;
			14'd2541: ff_rdata <= 8'h00;
			14'd2542: ff_rdata <= 8'h90;
			14'd2543: ff_rdata <= 8'h48;
			14'd2544: ff_rdata <= 8'h00;
			14'd2545: ff_rdata <= 8'h00;
			14'd2546: ff_rdata <= 8'h00;
			14'd2547: ff_rdata <= 8'h00;
			14'd2548: ff_rdata <= 8'h00;
			14'd2549: ff_rdata <= 8'h00;
			14'd2550: ff_rdata <= 8'h60;
			14'd2551: ff_rdata <= 8'h90;
			14'd2552: ff_rdata <= 8'h60;
			14'd2553: ff_rdata <= 8'h00;
			14'd2554: ff_rdata <= 8'h00;
			14'd2555: ff_rdata <= 8'h00;
			14'd2556: ff_rdata <= 8'h00;
			14'd2557: ff_rdata <= 8'h00;
			14'd2558: ff_rdata <= 8'h20;
			14'd2559: ff_rdata <= 8'hF8;
			14'd2560: ff_rdata <= 8'h20;
			14'd2561: ff_rdata <= 8'h4E;
			14'd2562: ff_rdata <= 8'h40;
			14'd2563: ff_rdata <= 8'h90;
			14'd2564: ff_rdata <= 8'h8E;
			14'd2565: ff_rdata <= 8'h00;
			14'd2566: ff_rdata <= 8'h10;
			14'd2567: ff_rdata <= 8'hFE;
			14'd2568: ff_rdata <= 8'h20;
			14'd2569: ff_rdata <= 8'h78;
			14'd2570: ff_rdata <= 8'h04;
			14'd2571: ff_rdata <= 8'h04;
			14'd2572: ff_rdata <= 8'h78;
			14'd2573: ff_rdata <= 8'h00;
			14'd2574: ff_rdata <= 8'h00;
			14'd2575: ff_rdata <= 8'hFC;
			14'd2576: ff_rdata <= 8'h02;
			14'd2577: ff_rdata <= 8'h02;
			14'd2578: ff_rdata <= 8'h02;
			14'd2579: ff_rdata <= 8'h04;
			14'd2580: ff_rdata <= 8'h18;
			14'd2581: ff_rdata <= 8'h00;
			14'd2582: ff_rdata <= 8'hFE;
			14'd2583: ff_rdata <= 8'h08;
			14'd2584: ff_rdata <= 8'h10;
			14'd2585: ff_rdata <= 8'h20;
			14'd2586: ff_rdata <= 8'h20;
			14'd2587: ff_rdata <= 8'h20;
			14'd2588: ff_rdata <= 8'h1C;
			14'd2589: ff_rdata <= 8'h00;
			14'd2590: ff_rdata <= 8'h20;
			14'd2591: ff_rdata <= 8'h24;
			14'd2592: ff_rdata <= 8'h38;
			14'd2593: ff_rdata <= 8'h60;
			14'd2594: ff_rdata <= 8'h80;
			14'd2595: ff_rdata <= 8'h80;
			14'd2596: ff_rdata <= 8'h7C;
			14'd2597: ff_rdata <= 8'h00;
			14'd2598: ff_rdata <= 8'h2C;
			14'd2599: ff_rdata <= 8'hF2;
			14'd2600: ff_rdata <= 8'h44;
			14'd2601: ff_rdata <= 8'h44;
			14'd2602: ff_rdata <= 8'h9C;
			14'd2603: ff_rdata <= 8'h26;
			14'd2604: ff_rdata <= 8'h1C;
			14'd2605: ff_rdata <= 8'h00;
			14'd2606: ff_rdata <= 8'h00;
			14'd2607: ff_rdata <= 8'h9E;
			14'd2608: ff_rdata <= 8'h80;
			14'd2609: ff_rdata <= 8'h80;
			14'd2610: ff_rdata <= 8'h80;
			14'd2611: ff_rdata <= 8'h90;
			14'd2612: ff_rdata <= 8'h4E;
			14'd2613: ff_rdata <= 8'h00;
			14'd2614: ff_rdata <= 8'h48;
			14'd2615: ff_rdata <= 8'h48;
			14'd2616: ff_rdata <= 8'h7C;
			14'd2617: ff_rdata <= 8'hD2;
			14'd2618: ff_rdata <= 8'hB6;
			14'd2619: ff_rdata <= 8'hAA;
			14'd2620: ff_rdata <= 8'h4C;
			14'd2621: ff_rdata <= 8'h00;
			14'd2622: ff_rdata <= 8'h40;
			14'd2623: ff_rdata <= 8'h4C;
			14'd2624: ff_rdata <= 8'hD2;
			14'd2625: ff_rdata <= 8'h62;
			14'd2626: ff_rdata <= 8'h4E;
			14'd2627: ff_rdata <= 8'hD2;
			14'd2628: ff_rdata <= 8'h4E;
			14'd2629: ff_rdata <= 8'h00;
			14'd2630: ff_rdata <= 8'h00;
			14'd2631: ff_rdata <= 8'h38;
			14'd2632: ff_rdata <= 8'h54;
			14'd2633: ff_rdata <= 8'h92;
			14'd2634: ff_rdata <= 8'hA2;
			14'd2635: ff_rdata <= 8'hA2;
			14'd2636: ff_rdata <= 8'h44;
			14'd2637: ff_rdata <= 8'h00;
			14'd2638: ff_rdata <= 8'h04;
			14'd2639: ff_rdata <= 8'h9E;
			14'd2640: ff_rdata <= 8'h84;
			14'd2641: ff_rdata <= 8'h84;
			14'd2642: ff_rdata <= 8'h8C;
			14'd2643: ff_rdata <= 8'h96;
			14'd2644: ff_rdata <= 8'h4C;
			14'd2645: ff_rdata <= 8'h00;
			14'd2646: ff_rdata <= 8'h10;
			14'd2647: ff_rdata <= 8'hE4;
			14'd2648: ff_rdata <= 8'h26;
			14'd2649: ff_rdata <= 8'h44;
			14'd2650: ff_rdata <= 8'h44;
			14'd2651: ff_rdata <= 8'h48;
			14'd2652: ff_rdata <= 8'h30;
			14'd2653: ff_rdata <= 8'h00;
			14'd2654: ff_rdata <= 8'h20;
			14'd2655: ff_rdata <= 8'h10;
			14'd2656: ff_rdata <= 8'h00;
			14'd2657: ff_rdata <= 8'h20;
			14'd2658: ff_rdata <= 8'h14;
			14'd2659: ff_rdata <= 8'h52;
			14'd2660: ff_rdata <= 8'hB2;
			14'd2661: ff_rdata <= 8'h00;
			14'd2662: ff_rdata <= 8'h00;
			14'd2663: ff_rdata <= 8'h00;
			14'd2664: ff_rdata <= 8'h20;
			14'd2665: ff_rdata <= 8'h50;
			14'd2666: ff_rdata <= 8'h88;
			14'd2667: ff_rdata <= 8'h04;
			14'd2668: ff_rdata <= 8'h02;
			14'd2669: ff_rdata <= 8'h00;
			14'd2670: ff_rdata <= 8'h1E;
			14'd2671: ff_rdata <= 8'h84;
			14'd2672: ff_rdata <= 8'h9E;
			14'd2673: ff_rdata <= 8'h84;
			14'd2674: ff_rdata <= 8'h8C;
			14'd2675: ff_rdata <= 8'h96;
			14'd2676: ff_rdata <= 8'h4C;
			14'd2677: ff_rdata <= 8'h00;
			14'd2678: ff_rdata <= 8'h10;
			14'd2679: ff_rdata <= 8'hFC;
			14'd2680: ff_rdata <= 8'h10;
			14'd2681: ff_rdata <= 8'hFC;
			14'd2682: ff_rdata <= 8'h70;
			14'd2683: ff_rdata <= 8'h98;
			14'd2684: ff_rdata <= 8'h74;
			14'd2685: ff_rdata <= 8'h00;
			14'd2686: ff_rdata <= 8'h70;
			14'd2687: ff_rdata <= 8'h10;
			14'd2688: ff_rdata <= 8'h14;
			14'd2689: ff_rdata <= 8'h7E;
			14'd2690: ff_rdata <= 8'hA4;
			14'd2691: ff_rdata <= 8'hA4;
			14'd2692: ff_rdata <= 8'h48;
			14'd2693: ff_rdata <= 8'h00;
			14'd2694: ff_rdata <= 8'h20;
			14'd2695: ff_rdata <= 8'hF4;
			14'd2696: ff_rdata <= 8'h22;
			14'd2697: ff_rdata <= 8'h60;
			14'd2698: ff_rdata <= 8'hA2;
			14'd2699: ff_rdata <= 8'h62;
			14'd2700: ff_rdata <= 8'h1C;
			14'd2701: ff_rdata <= 8'h00;
			14'd2702: ff_rdata <= 8'h48;
			14'd2703: ff_rdata <= 8'h48;
			14'd2704: ff_rdata <= 8'h7C;
			14'd2705: ff_rdata <= 8'hAA;
			14'd2706: ff_rdata <= 8'h92;
			14'd2707: ff_rdata <= 8'hA2;
			14'd2708: ff_rdata <= 8'h44;
			14'd2709: ff_rdata <= 8'h00;
			14'd2710: ff_rdata <= 8'h20;
			14'd2711: ff_rdata <= 8'hF8;
			14'd2712: ff_rdata <= 8'h20;
			14'd2713: ff_rdata <= 8'hF8;
			14'd2714: ff_rdata <= 8'h20;
			14'd2715: ff_rdata <= 8'h24;
			14'd2716: ff_rdata <= 8'h18;
			14'd2717: ff_rdata <= 8'h00;
			14'd2718: ff_rdata <= 8'h48;
			14'd2719: ff_rdata <= 8'h5C;
			14'd2720: ff_rdata <= 8'h6A;
			14'd2721: ff_rdata <= 8'hE2;
			14'd2722: ff_rdata <= 8'h24;
			14'd2723: ff_rdata <= 8'h10;
			14'd2724: ff_rdata <= 8'h10;
			14'd2725: ff_rdata <= 8'h00;
			14'd2726: ff_rdata <= 8'h10;
			14'd2727: ff_rdata <= 8'h9C;
			14'd2728: ff_rdata <= 8'hB2;
			14'd2729: ff_rdata <= 8'hD2;
			14'd2730: ff_rdata <= 8'h92;
			14'd2731: ff_rdata <= 8'h1C;
			14'd2732: ff_rdata <= 8'h20;
			14'd2733: ff_rdata <= 8'h00;
			14'd2734: ff_rdata <= 8'h10;
			14'd2735: ff_rdata <= 8'h1C;
			14'd2736: ff_rdata <= 8'h10;
			14'd2737: ff_rdata <= 8'h10;
			14'd2738: ff_rdata <= 8'h78;
			14'd2739: ff_rdata <= 8'h94;
			14'd2740: ff_rdata <= 8'h70;
			14'd2741: ff_rdata <= 8'h00;
			14'd2742: ff_rdata <= 8'h60;
			14'd2743: ff_rdata <= 8'h10;
			14'd2744: ff_rdata <= 8'h80;
			14'd2745: ff_rdata <= 8'hB8;
			14'd2746: ff_rdata <= 8'hC4;
			14'd2747: ff_rdata <= 8'h84;
			14'd2748: ff_rdata <= 8'h38;
			14'd2749: ff_rdata <= 8'h00;
			14'd2750: ff_rdata <= 8'h08;
			14'd2751: ff_rdata <= 8'h84;
			14'd2752: ff_rdata <= 8'h84;
			14'd2753: ff_rdata <= 8'h84;
			14'd2754: ff_rdata <= 8'h44;
			14'd2755: ff_rdata <= 8'h08;
			14'd2756: ff_rdata <= 8'h30;
			14'd2757: ff_rdata <= 8'h00;
			14'd2758: ff_rdata <= 8'h78;
			14'd2759: ff_rdata <= 8'h10;
			14'd2760: ff_rdata <= 8'h38;
			14'd2761: ff_rdata <= 8'h44;
			14'd2762: ff_rdata <= 8'hB4;
			14'd2763: ff_rdata <= 8'h4C;
			14'd2764: ff_rdata <= 8'h38;
			14'd2765: ff_rdata <= 8'h00;
			14'd2766: ff_rdata <= 8'h20;
			14'd2767: ff_rdata <= 8'h2C;
			14'd2768: ff_rdata <= 8'hF4;
			14'd2769: ff_rdata <= 8'h24;
			14'd2770: ff_rdata <= 8'h64;
			14'd2771: ff_rdata <= 8'hA4;
			14'd2772: ff_rdata <= 8'h26;
			14'd2773: ff_rdata <= 8'h00;
			14'd2774: ff_rdata <= 8'h78;
			14'd2775: ff_rdata <= 8'h10;
			14'd2776: ff_rdata <= 8'h20;
			14'd2777: ff_rdata <= 8'h78;
			14'd2778: ff_rdata <= 8'h84;
			14'd2779: ff_rdata <= 8'h04;
			14'd2780: ff_rdata <= 8'h38;
			14'd2781: ff_rdata <= 8'h00;
			14'd2782: ff_rdata <= 8'h40;
			14'd2783: ff_rdata <= 8'h40;
			14'd2784: ff_rdata <= 8'hDC;
			14'd2785: ff_rdata <= 8'h62;
			14'd2786: ff_rdata <= 8'h42;
			14'd2787: ff_rdata <= 8'hC2;
			14'd2788: ff_rdata <= 8'h44;
			14'd2789: ff_rdata <= 8'h00;
			14'd2790: ff_rdata <= 8'h10;
			14'd2791: ff_rdata <= 8'h10;
			14'd2792: ff_rdata <= 8'h20;
			14'd2793: ff_rdata <= 8'h20;
			14'd2794: ff_rdata <= 8'h60;
			14'd2795: ff_rdata <= 8'h52;
			14'd2796: ff_rdata <= 8'h8C;
			14'd2797: ff_rdata <= 8'h00;
			14'd2798: ff_rdata <= 8'h00;
			14'd2799: ff_rdata <= 8'h00;
			14'd2800: ff_rdata <= 8'h00;
			14'd2801: ff_rdata <= 8'h00;
			14'd2802: ff_rdata <= 8'h00;
			14'd2803: ff_rdata <= 8'h00;
			14'd2804: ff_rdata <= 8'h00;
			14'd2805: ff_rdata <= 8'h00;
			14'd2806: ff_rdata <= 8'hFF;
			14'd2807: ff_rdata <= 8'hFF;
			14'd2808: ff_rdata <= 8'hFF;
			14'd2809: ff_rdata <= 8'hFF;
			14'd2810: ff_rdata <= 8'hFF;
			14'd2811: ff_rdata <= 8'hFF;
			14'd2812: ff_rdata <= 8'hFF;
			14'd2813: ff_rdata <= 8'hFF;
			default: ff_rdata <= 8'd0;
			endcase
			ff_rdata_en <= 1'b1;
		end
		else begin
			ff_rdata <= 8'd0;
			ff_rdata_en <= 1'b0;
		end
	end

	assign rdata	= ff_rdata;
	assign rdata_en	= ff_rdata_en;
endmodule
