`define MODULE_NAME SSCPLL_Top
`define DEVICE_25
