// -----------------------------------------------------------------------------
//	ip_sdram_dummy2.v
//	Copyright (C)2024 Takayuki Hara (HRA!)
//	
//	 Permission is hereby granted, free of charge, to any person obtaining a 
//	copy of this software and associated documentation files (the "Software"), 
//	to deal in the Software without restriction, including without limitation 
//	the rights to use, copy, modify, merge, publish, distribute, sublicense, 
//	and/or sell copies of the Software, and to permit persons to whom the 
//	Software is furnished to do so, subject to the following conditions:
//	
//	The above copyright notice and this permission notice shall be included in 
//	all copies or substantial portions of the Software.
//	
//	The Software is provided "as is", without warranty of any kind, express or 
//	implied, including but not limited to the warranties of merchantability, 
//	fitness for a particular purpose and noninfringement. In no event shall the 
//	authors or copyright holders be liable for any claim, damages or other 
//	liability, whether in an action of contract, tort or otherwise, arising 
//	from, out of or in connection with the Software or the use or other dealings 
//	in the Software.
// -----------------------------------------------------------------------------
//	Description:
//		Debugger
// -----------------------------------------------------------------------------

module ip_sdram (
	input				n_reset			,
	input				clk				,
	input				clk_sdram		,
	input				rd_n			,
	input				wr_n			,
	output				busy			,
	input	[16:0]		address			,
	input	[7:0]		wdata			,
	output	[15:0]		rdata			,
	output				rdata_en		,
	output				O_sdram_clk		,
	output				O_sdram_cke		,
	output				O_sdram_cs_n	,
	output				O_sdram_ras_n	,
	output				O_sdram_cas_n	,
	output				O_sdram_wen_n	,
	inout	[31:0]		IO_sdram_dq		,
	output	[10:0]		O_sdram_addr	,
	output	[1:0]		O_sdram_ba		,
	output	[3:0]		O_sdram_dqm		
);
	reg		[ 7:0]	ff_dbi;

	assign O_sdram_clk		= 1'b0;
	assign O_sdram_cke		= 1'b0;
	assign O_sdram_cs_n		= 1'b0;
	assign O_sdram_ras_n	= 1'b0;
	assign O_sdram_cas_n	= 1'b0;
	assign O_sdram_wen_n	= 1'b0;
	assign IO_sdram_dq		= 32'hZ;
	assign O_sdram_addr		= 11'd0;
	assign O_sdram_ba		= 2'b00;
	assign O_sdram_dqm		= 4'b0000;

	assign busy				= 1'b0;
	assign rdata			= { ff_dbi, ff_dbi };
	assign rdata_en			= 1'b0;

	always @( posedge clk ) begin
		case( address[13:0] )
		14'h0000:	ff_dbi <= 8'h00;
		14'h0001:	ff_dbi <= 8'h00;
		14'h0002:	ff_dbi <= 8'h00;
		14'h0003:	ff_dbi <= 8'h00;
		14'h0004:	ff_dbi <= 8'h00;
		14'h0005:	ff_dbi <= 8'h00;
		14'h0006:	ff_dbi <= 8'h00;
		14'h0007:	ff_dbi <= 8'h00;
		14'h0008:	ff_dbi <= 8'h7e;
		14'h0009:	ff_dbi <= 8'h42;
		14'h000a:	ff_dbi <= 8'h7e;
		14'h000b:	ff_dbi <= 8'h42;
		14'h000c:	ff_dbi <= 8'h7e;
		14'h000d:	ff_dbi <= 8'h42;
		14'h000e:	ff_dbi <= 8'h82;
		14'h000f:	ff_dbi <= 8'h00;
		14'h0010:	ff_dbi <= 8'h10;
		14'h0011:	ff_dbi <= 8'h92;
		14'h0012:	ff_dbi <= 8'h54;
		14'h0013:	ff_dbi <= 8'h10;
		14'h0014:	ff_dbi <= 8'h28;
		14'h0015:	ff_dbi <= 8'h44;
		14'h0016:	ff_dbi <= 8'h82;
		14'h0017:	ff_dbi <= 8'h00;
		14'h0018:	ff_dbi <= 8'h12;
		14'h0019:	ff_dbi <= 8'h14;
		14'h001a:	ff_dbi <= 8'hf8;
		14'h001b:	ff_dbi <= 8'h14;
		14'h001c:	ff_dbi <= 8'h34;
		14'h001d:	ff_dbi <= 8'h52;
		14'h001e:	ff_dbi <= 8'h92;
		14'h001f:	ff_dbi <= 8'h00;
		14'h0020:	ff_dbi <= 8'h10;
		14'h0021:	ff_dbi <= 8'h10;
		14'h0022:	ff_dbi <= 8'hfe;
		14'h0023:	ff_dbi <= 8'h10;
		14'h0024:	ff_dbi <= 8'h38;
		14'h0025:	ff_dbi <= 8'h54;
		14'h0026:	ff_dbi <= 8'h92;
		14'h0027:	ff_dbi <= 8'h00;
		14'h0028:	ff_dbi <= 8'h10;
		14'h0029:	ff_dbi <= 8'h28;
		14'h002a:	ff_dbi <= 8'h7c;
		14'h002b:	ff_dbi <= 8'h92;
		14'h002c:	ff_dbi <= 8'h38;
		14'h002d:	ff_dbi <= 8'h54;
		14'h002e:	ff_dbi <= 8'hfe;
		14'h002f:	ff_dbi <= 8'h00;
		14'h0030:	ff_dbi <= 8'h10;
		14'h0031:	ff_dbi <= 8'h10;
		14'h0032:	ff_dbi <= 8'h10;
		14'h0033:	ff_dbi <= 8'h7c;
		14'h0034:	ff_dbi <= 8'h10;
		14'h0035:	ff_dbi <= 8'h10;
		14'h0036:	ff_dbi <= 8'hfe;
		14'h0037:	ff_dbi <= 8'h00;
		14'h0038:	ff_dbi <= 8'h7e;
		14'h0039:	ff_dbi <= 8'h42;
		14'h003a:	ff_dbi <= 8'h42;
		14'h003b:	ff_dbi <= 8'h7e;
		14'h003c:	ff_dbi <= 8'h42;
		14'h003d:	ff_dbi <= 8'h42;
		14'h003e:	ff_dbi <= 8'h7e;
		14'h003f:	ff_dbi <= 8'h00;
		14'h0040:	ff_dbi <= 8'h40;
		14'h0041:	ff_dbi <= 8'h7e;
		14'h0042:	ff_dbi <= 8'h48;
		14'h0043:	ff_dbi <= 8'h3c;
		14'h0044:	ff_dbi <= 8'h28;
		14'h0045:	ff_dbi <= 8'h7e;
		14'h0046:	ff_dbi <= 8'h08;
		14'h0047:	ff_dbi <= 8'h00;
		14'h0048:	ff_dbi <= 8'hfe;
		14'h0049:	ff_dbi <= 8'h92;
		14'h004a:	ff_dbi <= 8'h92;
		14'h004b:	ff_dbi <= 8'hfe;
		14'h004c:	ff_dbi <= 8'h82;
		14'h004d:	ff_dbi <= 8'h82;
		14'h004e:	ff_dbi <= 8'h86;
		14'h004f:	ff_dbi <= 8'h00;
		14'h0050:	ff_dbi <= 8'h04;
		14'h0051:	ff_dbi <= 8'hee;
		14'h0052:	ff_dbi <= 8'ha4;
		14'h0053:	ff_dbi <= 8'hef;
		14'h0054:	ff_dbi <= 8'ha2;
		14'h0055:	ff_dbi <= 8'hea;
		14'h0056:	ff_dbi <= 8'h06;
		14'h0057:	ff_dbi <= 8'h00;
		14'h0058:	ff_dbi <= 8'h28;
		14'h0059:	ff_dbi <= 8'h44;
		14'h005a:	ff_dbi <= 8'h82;
		14'h005b:	ff_dbi <= 8'h3c;
		14'h005c:	ff_dbi <= 8'h14;
		14'h005d:	ff_dbi <= 8'h24;
		14'h005e:	ff_dbi <= 8'h4c;
		14'h005f:	ff_dbi <= 8'h00;
		14'h0060:	ff_dbi <= 8'h28;
		14'h0061:	ff_dbi <= 8'hc8;
		14'h0062:	ff_dbi <= 8'h5c;
		14'h0063:	ff_dbi <= 8'hea;
		14'h0064:	ff_dbi <= 8'h6c;
		14'h0065:	ff_dbi <= 8'hc8;
		14'h0066:	ff_dbi <= 8'h50;
		14'h0067:	ff_dbi <= 8'h00;
		14'h0068:	ff_dbi <= 8'h7c;
		14'h0069:	ff_dbi <= 8'h20;
		14'h006a:	ff_dbi <= 8'h7c;
		14'h006b:	ff_dbi <= 8'h44;
		14'h006c:	ff_dbi <= 8'h7c;
		14'h006d:	ff_dbi <= 8'h44;
		14'h006e:	ff_dbi <= 8'h7c;
		14'h006f:	ff_dbi <= 8'h00;
		14'h0070:	ff_dbi <= 8'h0c;
		14'h0071:	ff_dbi <= 8'h70;
		14'h0072:	ff_dbi <= 8'h10;
		14'h0073:	ff_dbi <= 8'hfe;
		14'h0074:	ff_dbi <= 8'h10;
		14'h0075:	ff_dbi <= 8'h10;
		14'h0076:	ff_dbi <= 8'h10;
		14'h0077:	ff_dbi <= 8'h00;
		14'h0078:	ff_dbi <= 8'h7e;
		14'h0079:	ff_dbi <= 8'h10;
		14'h007a:	ff_dbi <= 8'h1e;
		14'h007b:	ff_dbi <= 8'h12;
		14'h007c:	ff_dbi <= 8'h22;
		14'h007d:	ff_dbi <= 8'h44;
		14'h007e:	ff_dbi <= 8'h08;
		14'h007f:	ff_dbi <= 8'h00;
		14'h0080:	ff_dbi <= 8'h00;
		14'h0081:	ff_dbi <= 8'h7c;
		14'h0082:	ff_dbi <= 8'h28;
		14'h0083:	ff_dbi <= 8'h28;
		14'h0084:	ff_dbi <= 8'h28;
		14'h0085:	ff_dbi <= 8'h4e;
		14'h0086:	ff_dbi <= 8'h00;
		14'h0087:	ff_dbi <= 8'h00;
		14'h0088:	ff_dbi <= 8'h10;
		14'h0089:	ff_dbi <= 8'h10;
		14'h008a:	ff_dbi <= 8'h10;
		14'h008b:	ff_dbi <= 8'hff;
		14'h008c:	ff_dbi <= 8'h00;
		14'h008d:	ff_dbi <= 8'h00;
		14'h008e:	ff_dbi <= 8'h00;
		14'h008f:	ff_dbi <= 8'h00;
		14'h0090:	ff_dbi <= 8'h00;
		14'h0091:	ff_dbi <= 8'h00;
		14'h0092:	ff_dbi <= 8'h00;
		14'h0093:	ff_dbi <= 8'hff;
		14'h0094:	ff_dbi <= 8'h10;
		14'h0095:	ff_dbi <= 8'h10;
		14'h0096:	ff_dbi <= 8'h10;
		14'h0097:	ff_dbi <= 8'h10;
		14'h0098:	ff_dbi <= 8'h10;
		14'h0099:	ff_dbi <= 8'h10;
		14'h009a:	ff_dbi <= 8'h10;
		14'h009b:	ff_dbi <= 8'hf0;
		14'h009c:	ff_dbi <= 8'h10;
		14'h009d:	ff_dbi <= 8'h10;
		14'h009e:	ff_dbi <= 8'h10;
		14'h009f:	ff_dbi <= 8'h10;
		14'h00a0:	ff_dbi <= 8'h10;
		14'h00a1:	ff_dbi <= 8'h10;
		14'h00a2:	ff_dbi <= 8'h10;
		14'h00a3:	ff_dbi <= 8'h1f;
		14'h00a4:	ff_dbi <= 8'h10;
		14'h00a5:	ff_dbi <= 8'h10;
		14'h00a6:	ff_dbi <= 8'h10;
		14'h00a7:	ff_dbi <= 8'h10;
		14'h00a8:	ff_dbi <= 8'h10;
		14'h00a9:	ff_dbi <= 8'h10;
		14'h00aa:	ff_dbi <= 8'h10;
		14'h00ab:	ff_dbi <= 8'hff;
		14'h00ac:	ff_dbi <= 8'h10;
		14'h00ad:	ff_dbi <= 8'h10;
		14'h00ae:	ff_dbi <= 8'h10;
		14'h00af:	ff_dbi <= 8'h10;
		14'h00b0:	ff_dbi <= 8'h10;
		14'h00b1:	ff_dbi <= 8'h10;
		14'h00b2:	ff_dbi <= 8'h10;
		14'h00b3:	ff_dbi <= 8'h10;
		14'h00b4:	ff_dbi <= 8'h10;
		14'h00b5:	ff_dbi <= 8'h10;
		14'h00b6:	ff_dbi <= 8'h10;
		14'h00b7:	ff_dbi <= 8'h10;
		14'h00b8:	ff_dbi <= 8'h00;
		14'h00b9:	ff_dbi <= 8'h00;
		14'h00ba:	ff_dbi <= 8'h00;
		14'h00bb:	ff_dbi <= 8'hff;
		14'h00bc:	ff_dbi <= 8'h00;
		14'h00bd:	ff_dbi <= 8'h00;
		14'h00be:	ff_dbi <= 8'h00;
		14'h00bf:	ff_dbi <= 8'h00;
		14'h00c0:	ff_dbi <= 8'h00;
		14'h00c1:	ff_dbi <= 8'h00;
		14'h00c2:	ff_dbi <= 8'h00;
		14'h00c3:	ff_dbi <= 8'h1f;
		14'h00c4:	ff_dbi <= 8'h10;
		14'h00c5:	ff_dbi <= 8'h10;
		14'h00c6:	ff_dbi <= 8'h10;
		14'h00c7:	ff_dbi <= 8'h10;
		14'h00c8:	ff_dbi <= 8'h00;
		14'h00c9:	ff_dbi <= 8'h00;
		14'h00ca:	ff_dbi <= 8'h00;
		14'h00cb:	ff_dbi <= 8'hf0;
		14'h00cc:	ff_dbi <= 8'h10;
		14'h00cd:	ff_dbi <= 8'h10;
		14'h00ce:	ff_dbi <= 8'h10;
		14'h00cf:	ff_dbi <= 8'h10;
		14'h00d0:	ff_dbi <= 8'h10;
		14'h00d1:	ff_dbi <= 8'h10;
		14'h00d2:	ff_dbi <= 8'h10;
		14'h00d3:	ff_dbi <= 8'h1f;
		14'h00d4:	ff_dbi <= 8'h00;
		14'h00d5:	ff_dbi <= 8'h00;
		14'h00d6:	ff_dbi <= 8'h00;
		14'h00d7:	ff_dbi <= 8'h00;
		14'h00d8:	ff_dbi <= 8'h10;
		14'h00d9:	ff_dbi <= 8'h10;
		14'h00da:	ff_dbi <= 8'h10;
		14'h00db:	ff_dbi <= 8'hf0;
		14'h00dc:	ff_dbi <= 8'h00;
		14'h00dd:	ff_dbi <= 8'h00;
		14'h00de:	ff_dbi <= 8'h00;
		14'h00df:	ff_dbi <= 8'h00;
		14'h00e0:	ff_dbi <= 8'h81;
		14'h00e1:	ff_dbi <= 8'h42;
		14'h00e2:	ff_dbi <= 8'h24;
		14'h00e3:	ff_dbi <= 8'h18;
		14'h00e4:	ff_dbi <= 8'h18;
		14'h00e5:	ff_dbi <= 8'h24;
		14'h00e6:	ff_dbi <= 8'h42;
		14'h00e7:	ff_dbi <= 8'h81;
		14'h00e8:	ff_dbi <= 8'h10;
		14'h00e9:	ff_dbi <= 8'h7c;
		14'h00ea:	ff_dbi <= 8'h10;
		14'h00eb:	ff_dbi <= 8'h10;
		14'h00ec:	ff_dbi <= 8'h28;
		14'h00ed:	ff_dbi <= 8'h44;
		14'h00ee:	ff_dbi <= 8'h82;
		14'h00ef:	ff_dbi <= 8'h00;
		14'h00f0:	ff_dbi <= 8'h10;
		14'h00f1:	ff_dbi <= 8'h10;
		14'h00f2:	ff_dbi <= 8'hfe;
		14'h00f3:	ff_dbi <= 8'h92;
		14'h00f4:	ff_dbi <= 8'hfe;
		14'h00f5:	ff_dbi <= 8'h10;
		14'h00f6:	ff_dbi <= 8'h10;
		14'h00f7:	ff_dbi <= 8'h00;
		14'h00f8:	ff_dbi <= 8'h10;
		14'h00f9:	ff_dbi <= 8'h10;
		14'h00fa:	ff_dbi <= 8'h54;
		14'h00fb:	ff_dbi <= 8'h54;
		14'h00fc:	ff_dbi <= 8'h92;
		14'h00fd:	ff_dbi <= 8'h10;
		14'h00fe:	ff_dbi <= 8'h30;
		14'h00ff:	ff_dbi <= 8'h00;
		14'h0100:	ff_dbi <= 8'h00;
		14'h0101:	ff_dbi <= 8'h00;
		14'h0102:	ff_dbi <= 8'h00;
		14'h0103:	ff_dbi <= 8'h00;
		14'h0104:	ff_dbi <= 8'h00;
		14'h0105:	ff_dbi <= 8'h00;
		14'h0106:	ff_dbi <= 8'h00;
		14'h0107:	ff_dbi <= 8'h00;
		14'h0108:	ff_dbi <= 8'h20;
		14'h0109:	ff_dbi <= 8'h20;
		14'h010a:	ff_dbi <= 8'h20;
		14'h010b:	ff_dbi <= 8'h20;
		14'h010c:	ff_dbi <= 8'h00;
		14'h010d:	ff_dbi <= 8'h00;
		14'h010e:	ff_dbi <= 8'h20;
		14'h010f:	ff_dbi <= 8'h00;
		14'h0110:	ff_dbi <= 8'h50;
		14'h0111:	ff_dbi <= 8'h50;
		14'h0112:	ff_dbi <= 8'h50;
		14'h0113:	ff_dbi <= 8'h00;
		14'h0114:	ff_dbi <= 8'h00;
		14'h0115:	ff_dbi <= 8'h00;
		14'h0116:	ff_dbi <= 8'h00;
		14'h0117:	ff_dbi <= 8'h00;
		14'h0118:	ff_dbi <= 8'h50;
		14'h0119:	ff_dbi <= 8'h50;
		14'h011a:	ff_dbi <= 8'hf8;
		14'h011b:	ff_dbi <= 8'h50;
		14'h011c:	ff_dbi <= 8'hf8;
		14'h011d:	ff_dbi <= 8'h50;
		14'h011e:	ff_dbi <= 8'h50;
		14'h011f:	ff_dbi <= 8'h00;
		14'h0120:	ff_dbi <= 8'h20;
		14'h0121:	ff_dbi <= 8'h78;
		14'h0122:	ff_dbi <= 8'ha0;
		14'h0123:	ff_dbi <= 8'h70;
		14'h0124:	ff_dbi <= 8'h28;
		14'h0125:	ff_dbi <= 8'hf0;
		14'h0126:	ff_dbi <= 8'h20;
		14'h0127:	ff_dbi <= 8'h00;
		14'h0128:	ff_dbi <= 8'hc0;
		14'h0129:	ff_dbi <= 8'hc8;
		14'h012a:	ff_dbi <= 8'h10;
		14'h012b:	ff_dbi <= 8'h20;
		14'h012c:	ff_dbi <= 8'h40;
		14'h012d:	ff_dbi <= 8'h98;
		14'h012e:	ff_dbi <= 8'h18;
		14'h012f:	ff_dbi <= 8'h00;
		14'h0130:	ff_dbi <= 8'h40;
		14'h0131:	ff_dbi <= 8'ha0;
		14'h0132:	ff_dbi <= 8'h40;
		14'h0133:	ff_dbi <= 8'ha8;
		14'h0134:	ff_dbi <= 8'h90;
		14'h0135:	ff_dbi <= 8'h98;
		14'h0136:	ff_dbi <= 8'h60;
		14'h0137:	ff_dbi <= 8'h00;
		14'h0138:	ff_dbi <= 8'h10;
		14'h0139:	ff_dbi <= 8'h20;
		14'h013a:	ff_dbi <= 8'h40;
		14'h013b:	ff_dbi <= 8'h00;
		14'h013c:	ff_dbi <= 8'h00;
		14'h013d:	ff_dbi <= 8'h00;
		14'h013e:	ff_dbi <= 8'h00;
		14'h013f:	ff_dbi <= 8'h00;
		14'h0140:	ff_dbi <= 8'h10;
		14'h0141:	ff_dbi <= 8'h20;
		14'h0142:	ff_dbi <= 8'h40;
		14'h0143:	ff_dbi <= 8'h40;
		14'h0144:	ff_dbi <= 8'h40;
		14'h0145:	ff_dbi <= 8'h20;
		14'h0146:	ff_dbi <= 8'h10;
		14'h0147:	ff_dbi <= 8'h00;
		14'h0148:	ff_dbi <= 8'h40;
		14'h0149:	ff_dbi <= 8'h20;
		14'h014a:	ff_dbi <= 8'h10;
		14'h014b:	ff_dbi <= 8'h10;
		14'h014c:	ff_dbi <= 8'h10;
		14'h014d:	ff_dbi <= 8'h20;
		14'h014e:	ff_dbi <= 8'h40;
		14'h014f:	ff_dbi <= 8'h00;
		14'h0150:	ff_dbi <= 8'h20;
		14'h0151:	ff_dbi <= 8'ha8;
		14'h0152:	ff_dbi <= 8'h70;
		14'h0153:	ff_dbi <= 8'h20;
		14'h0154:	ff_dbi <= 8'h70;
		14'h0155:	ff_dbi <= 8'ha8;
		14'h0156:	ff_dbi <= 8'h20;
		14'h0157:	ff_dbi <= 8'h00;
		14'h0158:	ff_dbi <= 8'h00;
		14'h0159:	ff_dbi <= 8'h20;
		14'h015a:	ff_dbi <= 8'h20;
		14'h015b:	ff_dbi <= 8'hf8;
		14'h015c:	ff_dbi <= 8'h20;
		14'h015d:	ff_dbi <= 8'h20;
		14'h015e:	ff_dbi <= 8'h00;
		14'h015f:	ff_dbi <= 8'h00;
		14'h0160:	ff_dbi <= 8'h00;
		14'h0161:	ff_dbi <= 8'h00;
		14'h0162:	ff_dbi <= 8'h00;
		14'h0163:	ff_dbi <= 8'h00;
		14'h0164:	ff_dbi <= 8'h00;
		14'h0165:	ff_dbi <= 8'h20;
		14'h0166:	ff_dbi <= 8'h20;
		14'h0167:	ff_dbi <= 8'h40;
		14'h0168:	ff_dbi <= 8'h00;
		14'h0169:	ff_dbi <= 8'h00;
		14'h016a:	ff_dbi <= 8'h00;
		14'h016b:	ff_dbi <= 8'h78;
		14'h016c:	ff_dbi <= 8'h00;
		14'h016d:	ff_dbi <= 8'h00;
		14'h016e:	ff_dbi <= 8'h00;
		14'h016f:	ff_dbi <= 8'h00;
		14'h0170:	ff_dbi <= 8'h00;
		14'h0171:	ff_dbi <= 8'h00;
		14'h0172:	ff_dbi <= 8'h00;
		14'h0173:	ff_dbi <= 8'h00;
		14'h0174:	ff_dbi <= 8'h00;
		14'h0175:	ff_dbi <= 8'h60;
		14'h0176:	ff_dbi <= 8'h60;
		14'h0177:	ff_dbi <= 8'h00;
		14'h0178:	ff_dbi <= 8'h00;
		14'h0179:	ff_dbi <= 8'h00;
		14'h017a:	ff_dbi <= 8'h08;
		14'h017b:	ff_dbi <= 8'h10;
		14'h017c:	ff_dbi <= 8'h20;
		14'h017d:	ff_dbi <= 8'h40;
		14'h017e:	ff_dbi <= 8'h80;
		14'h017f:	ff_dbi <= 8'h00;
		14'h0180:	ff_dbi <= 8'h70;
		14'h0181:	ff_dbi <= 8'h88;
		14'h0182:	ff_dbi <= 8'h98;
		14'h0183:	ff_dbi <= 8'ha8;
		14'h0184:	ff_dbi <= 8'hc8;
		14'h0185:	ff_dbi <= 8'h88;
		14'h0186:	ff_dbi <= 8'h70;
		14'h0187:	ff_dbi <= 8'h00;
		14'h0188:	ff_dbi <= 8'h20;
		14'h0189:	ff_dbi <= 8'h60;
		14'h018a:	ff_dbi <= 8'ha0;
		14'h018b:	ff_dbi <= 8'h20;
		14'h018c:	ff_dbi <= 8'h20;
		14'h018d:	ff_dbi <= 8'h20;
		14'h018e:	ff_dbi <= 8'hf8;
		14'h018f:	ff_dbi <= 8'h00;
		14'h0190:	ff_dbi <= 8'h70;
		14'h0191:	ff_dbi <= 8'h88;
		14'h0192:	ff_dbi <= 8'h08;
		14'h0193:	ff_dbi <= 8'h10;
		14'h0194:	ff_dbi <= 8'h60;
		14'h0195:	ff_dbi <= 8'h80;
		14'h0196:	ff_dbi <= 8'hf8;
		14'h0197:	ff_dbi <= 8'h00;
		14'h0198:	ff_dbi <= 8'h70;
		14'h0199:	ff_dbi <= 8'h88;
		14'h019a:	ff_dbi <= 8'h08;
		14'h019b:	ff_dbi <= 8'h30;
		14'h019c:	ff_dbi <= 8'h08;
		14'h019d:	ff_dbi <= 8'h88;
		14'h019e:	ff_dbi <= 8'h70;
		14'h019f:	ff_dbi <= 8'h00;
		14'h01a0:	ff_dbi <= 8'h10;
		14'h01a1:	ff_dbi <= 8'h30;
		14'h01a2:	ff_dbi <= 8'h50;
		14'h01a3:	ff_dbi <= 8'h90;
		14'h01a4:	ff_dbi <= 8'hf8;
		14'h01a5:	ff_dbi <= 8'h10;
		14'h01a6:	ff_dbi <= 8'h10;
		14'h01a7:	ff_dbi <= 8'h00;
		14'h01a8:	ff_dbi <= 8'hf8;
		14'h01a9:	ff_dbi <= 8'h80;
		14'h01aa:	ff_dbi <= 8'he0;
		14'h01ab:	ff_dbi <= 8'h10;
		14'h01ac:	ff_dbi <= 8'h08;
		14'h01ad:	ff_dbi <= 8'h10;
		14'h01ae:	ff_dbi <= 8'he0;
		14'h01af:	ff_dbi <= 8'h00;
		14'h01b0:	ff_dbi <= 8'h30;
		14'h01b1:	ff_dbi <= 8'h40;
		14'h01b2:	ff_dbi <= 8'h80;
		14'h01b3:	ff_dbi <= 8'hf0;
		14'h01b4:	ff_dbi <= 8'h88;
		14'h01b5:	ff_dbi <= 8'h88;
		14'h01b6:	ff_dbi <= 8'h70;
		14'h01b7:	ff_dbi <= 8'h00;
		14'h01b8:	ff_dbi <= 8'hf8;
		14'h01b9:	ff_dbi <= 8'h88;
		14'h01ba:	ff_dbi <= 8'h10;
		14'h01bb:	ff_dbi <= 8'h20;
		14'h01bc:	ff_dbi <= 8'h20;
		14'h01bd:	ff_dbi <= 8'h20;
		14'h01be:	ff_dbi <= 8'h20;
		14'h01bf:	ff_dbi <= 8'h00;
		14'h01c0:	ff_dbi <= 8'h70;
		14'h01c1:	ff_dbi <= 8'h88;
		14'h01c2:	ff_dbi <= 8'h88;
		14'h01c3:	ff_dbi <= 8'h70;
		14'h01c4:	ff_dbi <= 8'h88;
		14'h01c5:	ff_dbi <= 8'h88;
		14'h01c6:	ff_dbi <= 8'h70;
		14'h01c7:	ff_dbi <= 8'h00;
		14'h01c8:	ff_dbi <= 8'h70;
		14'h01c9:	ff_dbi <= 8'h88;
		14'h01ca:	ff_dbi <= 8'h88;
		14'h01cb:	ff_dbi <= 8'h78;
		14'h01cc:	ff_dbi <= 8'h08;
		14'h01cd:	ff_dbi <= 8'h10;
		14'h01ce:	ff_dbi <= 8'h60;
		14'h01cf:	ff_dbi <= 8'h00;
		14'h01d0:	ff_dbi <= 8'h00;
		14'h01d1:	ff_dbi <= 8'h00;
		14'h01d2:	ff_dbi <= 8'h20;
		14'h01d3:	ff_dbi <= 8'h00;
		14'h01d4:	ff_dbi <= 8'h00;
		14'h01d5:	ff_dbi <= 8'h20;
		14'h01d6:	ff_dbi <= 8'h00;
		14'h01d7:	ff_dbi <= 8'h00;
		14'h01d8:	ff_dbi <= 8'h00;
		14'h01d9:	ff_dbi <= 8'h00;
		14'h01da:	ff_dbi <= 8'h20;
		14'h01db:	ff_dbi <= 8'h00;
		14'h01dc:	ff_dbi <= 8'h00;
		14'h01dd:	ff_dbi <= 8'h20;
		14'h01de:	ff_dbi <= 8'h20;
		14'h01df:	ff_dbi <= 8'h40;
		14'h01e0:	ff_dbi <= 8'h18;
		14'h01e1:	ff_dbi <= 8'h30;
		14'h01e2:	ff_dbi <= 8'h60;
		14'h01e3:	ff_dbi <= 8'hc0;
		14'h01e4:	ff_dbi <= 8'h60;
		14'h01e5:	ff_dbi <= 8'h30;
		14'h01e6:	ff_dbi <= 8'h18;
		14'h01e7:	ff_dbi <= 8'h00;
		14'h01e8:	ff_dbi <= 8'h00;
		14'h01e9:	ff_dbi <= 8'h00;
		14'h01ea:	ff_dbi <= 8'hf8;
		14'h01eb:	ff_dbi <= 8'h00;
		14'h01ec:	ff_dbi <= 8'hf8;
		14'h01ed:	ff_dbi <= 8'h00;
		14'h01ee:	ff_dbi <= 8'h00;
		14'h01ef:	ff_dbi <= 8'h00;
		14'h01f0:	ff_dbi <= 8'hc0;
		14'h01f1:	ff_dbi <= 8'h60;
		14'h01f2:	ff_dbi <= 8'h30;
		14'h01f3:	ff_dbi <= 8'h18;
		14'h01f4:	ff_dbi <= 8'h30;
		14'h01f5:	ff_dbi <= 8'h60;
		14'h01f6:	ff_dbi <= 8'hc0;
		14'h01f7:	ff_dbi <= 8'h00;
		14'h01f8:	ff_dbi <= 8'h70;
		14'h01f9:	ff_dbi <= 8'h88;
		14'h01fa:	ff_dbi <= 8'h08;
		14'h01fb:	ff_dbi <= 8'h10;
		14'h01fc:	ff_dbi <= 8'h20;
		14'h01fd:	ff_dbi <= 8'h00;
		14'h01fe:	ff_dbi <= 8'h20;
		14'h01ff:	ff_dbi <= 8'h00;
		14'h0200:	ff_dbi <= 8'h70;
		14'h0201:	ff_dbi <= 8'h88;
		14'h0202:	ff_dbi <= 8'h08;
		14'h0203:	ff_dbi <= 8'h68;
		14'h0204:	ff_dbi <= 8'ha8;
		14'h0205:	ff_dbi <= 8'ha8;
		14'h0206:	ff_dbi <= 8'h70;
		14'h0207:	ff_dbi <= 8'h00;
		14'h0208:	ff_dbi <= 8'h20;
		14'h0209:	ff_dbi <= 8'h50;
		14'h020a:	ff_dbi <= 8'h88;
		14'h020b:	ff_dbi <= 8'h88;
		14'h020c:	ff_dbi <= 8'hf8;
		14'h020d:	ff_dbi <= 8'h88;
		14'h020e:	ff_dbi <= 8'h88;
		14'h020f:	ff_dbi <= 8'h00;
		14'h0210:	ff_dbi <= 8'hf0;
		14'h0211:	ff_dbi <= 8'h48;
		14'h0212:	ff_dbi <= 8'h48;
		14'h0213:	ff_dbi <= 8'h70;
		14'h0214:	ff_dbi <= 8'h48;
		14'h0215:	ff_dbi <= 8'h48;
		14'h0216:	ff_dbi <= 8'hf0;
		14'h0217:	ff_dbi <= 8'h00;
		14'h0218:	ff_dbi <= 8'h30;
		14'h0219:	ff_dbi <= 8'h48;
		14'h021a:	ff_dbi <= 8'h80;
		14'h021b:	ff_dbi <= 8'h80;
		14'h021c:	ff_dbi <= 8'h80;
		14'h021d:	ff_dbi <= 8'h48;
		14'h021e:	ff_dbi <= 8'h30;
		14'h021f:	ff_dbi <= 8'h00;
		14'h0220:	ff_dbi <= 8'he0;
		14'h0221:	ff_dbi <= 8'h50;
		14'h0222:	ff_dbi <= 8'h48;
		14'h0223:	ff_dbi <= 8'h48;
		14'h0224:	ff_dbi <= 8'h48;
		14'h0225:	ff_dbi <= 8'h50;
		14'h0226:	ff_dbi <= 8'he0;
		14'h0227:	ff_dbi <= 8'h00;
		14'h0228:	ff_dbi <= 8'hf8;
		14'h0229:	ff_dbi <= 8'h80;
		14'h022a:	ff_dbi <= 8'h80;
		14'h022b:	ff_dbi <= 8'hf0;
		14'h022c:	ff_dbi <= 8'h80;
		14'h022d:	ff_dbi <= 8'h80;
		14'h022e:	ff_dbi <= 8'hf8;
		14'h022f:	ff_dbi <= 8'h00;
		14'h0230:	ff_dbi <= 8'hf8;
		14'h0231:	ff_dbi <= 8'h80;
		14'h0232:	ff_dbi <= 8'h80;
		14'h0233:	ff_dbi <= 8'hf0;
		14'h0234:	ff_dbi <= 8'h80;
		14'h0235:	ff_dbi <= 8'h80;
		14'h0236:	ff_dbi <= 8'h80;
		14'h0237:	ff_dbi <= 8'h00;
		14'h0238:	ff_dbi <= 8'h70;
		14'h0239:	ff_dbi <= 8'h88;
		14'h023a:	ff_dbi <= 8'h80;
		14'h023b:	ff_dbi <= 8'hb8;
		14'h023c:	ff_dbi <= 8'h88;
		14'h023d:	ff_dbi <= 8'h88;
		14'h023e:	ff_dbi <= 8'h70;
		14'h023f:	ff_dbi <= 8'h00;
		14'h0240:	ff_dbi <= 8'h88;
		14'h0241:	ff_dbi <= 8'h88;
		14'h0242:	ff_dbi <= 8'h88;
		14'h0243:	ff_dbi <= 8'hf8;
		14'h0244:	ff_dbi <= 8'h88;
		14'h0245:	ff_dbi <= 8'h88;
		14'h0246:	ff_dbi <= 8'h88;
		14'h0247:	ff_dbi <= 8'h00;
		14'h0248:	ff_dbi <= 8'h70;
		14'h0249:	ff_dbi <= 8'h20;
		14'h024a:	ff_dbi <= 8'h20;
		14'h024b:	ff_dbi <= 8'h20;
		14'h024c:	ff_dbi <= 8'h20;
		14'h024d:	ff_dbi <= 8'h20;
		14'h024e:	ff_dbi <= 8'h70;
		14'h024f:	ff_dbi <= 8'h00;
		14'h0250:	ff_dbi <= 8'h38;
		14'h0251:	ff_dbi <= 8'h10;
		14'h0252:	ff_dbi <= 8'h10;
		14'h0253:	ff_dbi <= 8'h10;
		14'h0254:	ff_dbi <= 8'h90;
		14'h0255:	ff_dbi <= 8'h90;
		14'h0256:	ff_dbi <= 8'h60;
		14'h0257:	ff_dbi <= 8'h00;
		14'h0258:	ff_dbi <= 8'h88;
		14'h0259:	ff_dbi <= 8'h90;
		14'h025a:	ff_dbi <= 8'ha0;
		14'h025b:	ff_dbi <= 8'hc0;
		14'h025c:	ff_dbi <= 8'ha0;
		14'h025d:	ff_dbi <= 8'h90;
		14'h025e:	ff_dbi <= 8'h88;
		14'h025f:	ff_dbi <= 8'h00;
		14'h0260:	ff_dbi <= 8'h80;
		14'h0261:	ff_dbi <= 8'h80;
		14'h0262:	ff_dbi <= 8'h80;
		14'h0263:	ff_dbi <= 8'h80;
		14'h0264:	ff_dbi <= 8'h80;
		14'h0265:	ff_dbi <= 8'h80;
		14'h0266:	ff_dbi <= 8'hf8;
		14'h0267:	ff_dbi <= 8'h00;
		14'h0268:	ff_dbi <= 8'h88;
		14'h0269:	ff_dbi <= 8'hd8;
		14'h026a:	ff_dbi <= 8'ha8;
		14'h026b:	ff_dbi <= 8'ha8;
		14'h026c:	ff_dbi <= 8'h88;
		14'h026d:	ff_dbi <= 8'h88;
		14'h026e:	ff_dbi <= 8'h88;
		14'h026f:	ff_dbi <= 8'h00;
		14'h0270:	ff_dbi <= 8'h88;
		14'h0271:	ff_dbi <= 8'hc8;
		14'h0272:	ff_dbi <= 8'hc8;
		14'h0273:	ff_dbi <= 8'ha8;
		14'h0274:	ff_dbi <= 8'h98;
		14'h0275:	ff_dbi <= 8'h98;
		14'h0276:	ff_dbi <= 8'h88;
		14'h0277:	ff_dbi <= 8'h00;
		14'h0278:	ff_dbi <= 8'h70;
		14'h0279:	ff_dbi <= 8'h88;
		14'h027a:	ff_dbi <= 8'h88;
		14'h027b:	ff_dbi <= 8'h88;
		14'h027c:	ff_dbi <= 8'h88;
		14'h027d:	ff_dbi <= 8'h88;
		14'h027e:	ff_dbi <= 8'h70;
		14'h027f:	ff_dbi <= 8'h00;
		14'h0280:	ff_dbi <= 8'hf0;
		14'h0281:	ff_dbi <= 8'h88;
		14'h0282:	ff_dbi <= 8'h88;
		14'h0283:	ff_dbi <= 8'hf0;
		14'h0284:	ff_dbi <= 8'h80;
		14'h0285:	ff_dbi <= 8'h80;
		14'h0286:	ff_dbi <= 8'h80;
		14'h0287:	ff_dbi <= 8'h00;
		14'h0288:	ff_dbi <= 8'h70;
		14'h0289:	ff_dbi <= 8'h88;
		14'h028a:	ff_dbi <= 8'h88;
		14'h028b:	ff_dbi <= 8'h88;
		14'h028c:	ff_dbi <= 8'ha8;
		14'h028d:	ff_dbi <= 8'h90;
		14'h028e:	ff_dbi <= 8'h68;
		14'h028f:	ff_dbi <= 8'h00;
		14'h0290:	ff_dbi <= 8'hf0;
		14'h0291:	ff_dbi <= 8'h88;
		14'h0292:	ff_dbi <= 8'h88;
		14'h0293:	ff_dbi <= 8'hf0;
		14'h0294:	ff_dbi <= 8'ha0;
		14'h0295:	ff_dbi <= 8'h90;
		14'h0296:	ff_dbi <= 8'h88;
		14'h0297:	ff_dbi <= 8'h00;
		14'h0298:	ff_dbi <= 8'h70;
		14'h0299:	ff_dbi <= 8'h88;
		14'h029a:	ff_dbi <= 8'h80;
		14'h029b:	ff_dbi <= 8'h70;
		14'h029c:	ff_dbi <= 8'h08;
		14'h029d:	ff_dbi <= 8'h88;
		14'h029e:	ff_dbi <= 8'h70;
		14'h029f:	ff_dbi <= 8'h00;
		14'h02a0:	ff_dbi <= 8'hf8;
		14'h02a1:	ff_dbi <= 8'h20;
		14'h02a2:	ff_dbi <= 8'h20;
		14'h02a3:	ff_dbi <= 8'h20;
		14'h02a4:	ff_dbi <= 8'h20;
		14'h02a5:	ff_dbi <= 8'h20;
		14'h02a6:	ff_dbi <= 8'h20;
		14'h02a7:	ff_dbi <= 8'h00;
		14'h02a8:	ff_dbi <= 8'h88;
		14'h02a9:	ff_dbi <= 8'h88;
		14'h02aa:	ff_dbi <= 8'h88;
		14'h02ab:	ff_dbi <= 8'h88;
		14'h02ac:	ff_dbi <= 8'h88;
		14'h02ad:	ff_dbi <= 8'h88;
		14'h02ae:	ff_dbi <= 8'h70;
		14'h02af:	ff_dbi <= 8'h00;
		14'h02b0:	ff_dbi <= 8'h88;
		14'h02b1:	ff_dbi <= 8'h88;
		14'h02b2:	ff_dbi <= 8'h88;
		14'h02b3:	ff_dbi <= 8'h88;
		14'h02b4:	ff_dbi <= 8'h50;
		14'h02b5:	ff_dbi <= 8'h50;
		14'h02b6:	ff_dbi <= 8'h20;
		14'h02b7:	ff_dbi <= 8'h00;
		14'h02b8:	ff_dbi <= 8'h88;
		14'h02b9:	ff_dbi <= 8'h88;
		14'h02ba:	ff_dbi <= 8'h88;
		14'h02bb:	ff_dbi <= 8'ha8;
		14'h02bc:	ff_dbi <= 8'ha8;
		14'h02bd:	ff_dbi <= 8'hd8;
		14'h02be:	ff_dbi <= 8'h88;
		14'h02bf:	ff_dbi <= 8'h00;
		14'h02c0:	ff_dbi <= 8'h88;
		14'h02c1:	ff_dbi <= 8'h88;
		14'h02c2:	ff_dbi <= 8'h50;
		14'h02c3:	ff_dbi <= 8'h20;
		14'h02c4:	ff_dbi <= 8'h50;
		14'h02c5:	ff_dbi <= 8'h88;
		14'h02c6:	ff_dbi <= 8'h88;
		14'h02c7:	ff_dbi <= 8'h00;
		14'h02c8:	ff_dbi <= 8'h88;
		14'h02c9:	ff_dbi <= 8'h88;
		14'h02ca:	ff_dbi <= 8'h88;
		14'h02cb:	ff_dbi <= 8'h70;
		14'h02cc:	ff_dbi <= 8'h20;
		14'h02cd:	ff_dbi <= 8'h20;
		14'h02ce:	ff_dbi <= 8'h20;
		14'h02cf:	ff_dbi <= 8'h00;
		14'h02d0:	ff_dbi <= 8'hf8;
		14'h02d1:	ff_dbi <= 8'h08;
		14'h02d2:	ff_dbi <= 8'h10;
		14'h02d3:	ff_dbi <= 8'h20;
		14'h02d4:	ff_dbi <= 8'h40;
		14'h02d5:	ff_dbi <= 8'h80;
		14'h02d6:	ff_dbi <= 8'hf8;
		14'h02d7:	ff_dbi <= 8'h00;
		14'h02d8:	ff_dbi <= 8'h70;
		14'h02d9:	ff_dbi <= 8'h40;
		14'h02da:	ff_dbi <= 8'h40;
		14'h02db:	ff_dbi <= 8'h40;
		14'h02dc:	ff_dbi <= 8'h40;
		14'h02dd:	ff_dbi <= 8'h40;
		14'h02de:	ff_dbi <= 8'h70;
		14'h02df:	ff_dbi <= 8'h00;
		14'h02e0:	ff_dbi <= 8'h88;
		14'h02e1:	ff_dbi <= 8'h50;
		14'h02e2:	ff_dbi <= 8'h20;
		14'h02e3:	ff_dbi <= 8'h70;
		14'h02e4:	ff_dbi <= 8'h20;
		14'h02e5:	ff_dbi <= 8'h70;
		14'h02e6:	ff_dbi <= 8'h20;
		14'h02e7:	ff_dbi <= 8'h00;
		14'h02e8:	ff_dbi <= 8'h70;
		14'h02e9:	ff_dbi <= 8'h10;
		14'h02ea:	ff_dbi <= 8'h10;
		14'h02eb:	ff_dbi <= 8'h10;
		14'h02ec:	ff_dbi <= 8'h10;
		14'h02ed:	ff_dbi <= 8'h10;
		14'h02ee:	ff_dbi <= 8'h70;
		14'h02ef:	ff_dbi <= 8'h00;
		14'h02f0:	ff_dbi <= 8'h20;
		14'h02f1:	ff_dbi <= 8'h50;
		14'h02f2:	ff_dbi <= 8'h88;
		14'h02f3:	ff_dbi <= 8'h00;
		14'h02f4:	ff_dbi <= 8'h00;
		14'h02f5:	ff_dbi <= 8'h00;
		14'h02f6:	ff_dbi <= 8'h00;
		14'h02f7:	ff_dbi <= 8'h00;
		14'h02f8:	ff_dbi <= 8'h00;
		14'h02f9:	ff_dbi <= 8'h00;
		14'h02fa:	ff_dbi <= 8'h00;
		14'h02fb:	ff_dbi <= 8'h00;
		14'h02fc:	ff_dbi <= 8'h00;
		14'h02fd:	ff_dbi <= 8'h00;
		14'h02fe:	ff_dbi <= 8'hf8;
		14'h02ff:	ff_dbi <= 8'h00;
		14'h0300:	ff_dbi <= 8'h40;
		14'h0301:	ff_dbi <= 8'h20;
		14'h0302:	ff_dbi <= 8'h10;
		14'h0303:	ff_dbi <= 8'h00;
		14'h0304:	ff_dbi <= 8'h00;
		14'h0305:	ff_dbi <= 8'h00;
		14'h0306:	ff_dbi <= 8'h00;
		14'h0307:	ff_dbi <= 8'h00;
		14'h0308:	ff_dbi <= 8'h00;
		14'h0309:	ff_dbi <= 8'h00;
		14'h030a:	ff_dbi <= 8'h70;
		14'h030b:	ff_dbi <= 8'h08;
		14'h030c:	ff_dbi <= 8'h78;
		14'h030d:	ff_dbi <= 8'h88;
		14'h030e:	ff_dbi <= 8'h78;
		14'h030f:	ff_dbi <= 8'h00;
		14'h0310:	ff_dbi <= 8'h80;
		14'h0311:	ff_dbi <= 8'h80;
		14'h0312:	ff_dbi <= 8'hb0;
		14'h0313:	ff_dbi <= 8'hc8;
		14'h0314:	ff_dbi <= 8'h88;
		14'h0315:	ff_dbi <= 8'hc8;
		14'h0316:	ff_dbi <= 8'hb0;
		14'h0317:	ff_dbi <= 8'h00;
		14'h0318:	ff_dbi <= 8'h00;
		14'h0319:	ff_dbi <= 8'h00;
		14'h031a:	ff_dbi <= 8'h70;
		14'h031b:	ff_dbi <= 8'h88;
		14'h031c:	ff_dbi <= 8'h80;
		14'h031d:	ff_dbi <= 8'h88;
		14'h031e:	ff_dbi <= 8'h70;
		14'h031f:	ff_dbi <= 8'h00;
		14'h0320:	ff_dbi <= 8'h08;
		14'h0321:	ff_dbi <= 8'h08;
		14'h0322:	ff_dbi <= 8'h68;
		14'h0323:	ff_dbi <= 8'h98;
		14'h0324:	ff_dbi <= 8'h88;
		14'h0325:	ff_dbi <= 8'h98;
		14'h0326:	ff_dbi <= 8'h68;
		14'h0327:	ff_dbi <= 8'h00;
		14'h0328:	ff_dbi <= 8'h00;
		14'h0329:	ff_dbi <= 8'h00;
		14'h032a:	ff_dbi <= 8'h70;
		14'h032b:	ff_dbi <= 8'h88;
		14'h032c:	ff_dbi <= 8'hf8;
		14'h032d:	ff_dbi <= 8'h80;
		14'h032e:	ff_dbi <= 8'h70;
		14'h032f:	ff_dbi <= 8'h00;
		14'h0330:	ff_dbi <= 8'h10;
		14'h0331:	ff_dbi <= 8'h28;
		14'h0332:	ff_dbi <= 8'h20;
		14'h0333:	ff_dbi <= 8'hf8;
		14'h0334:	ff_dbi <= 8'h20;
		14'h0335:	ff_dbi <= 8'h20;
		14'h0336:	ff_dbi <= 8'h20;
		14'h0337:	ff_dbi <= 8'h00;
		14'h0338:	ff_dbi <= 8'h00;
		14'h0339:	ff_dbi <= 8'h00;
		14'h033a:	ff_dbi <= 8'h68;
		14'h033b:	ff_dbi <= 8'h98;
		14'h033c:	ff_dbi <= 8'h98;
		14'h033d:	ff_dbi <= 8'h68;
		14'h033e:	ff_dbi <= 8'h08;
		14'h033f:	ff_dbi <= 8'h70;
		14'h0340:	ff_dbi <= 8'h80;
		14'h0341:	ff_dbi <= 8'h80;
		14'h0342:	ff_dbi <= 8'hf0;
		14'h0343:	ff_dbi <= 8'h88;
		14'h0344:	ff_dbi <= 8'h88;
		14'h0345:	ff_dbi <= 8'h88;
		14'h0346:	ff_dbi <= 8'h88;
		14'h0347:	ff_dbi <= 8'h00;
		14'h0348:	ff_dbi <= 8'h20;
		14'h0349:	ff_dbi <= 8'h00;
		14'h034a:	ff_dbi <= 8'h60;
		14'h034b:	ff_dbi <= 8'h20;
		14'h034c:	ff_dbi <= 8'h20;
		14'h034d:	ff_dbi <= 8'h20;
		14'h034e:	ff_dbi <= 8'h70;
		14'h034f:	ff_dbi <= 8'h00;
		14'h0350:	ff_dbi <= 8'h10;
		14'h0351:	ff_dbi <= 8'h00;
		14'h0352:	ff_dbi <= 8'h30;
		14'h0353:	ff_dbi <= 8'h10;
		14'h0354:	ff_dbi <= 8'h10;
		14'h0355:	ff_dbi <= 8'h10;
		14'h0356:	ff_dbi <= 8'h90;
		14'h0357:	ff_dbi <= 8'h60;
		14'h0358:	ff_dbi <= 8'h40;
		14'h0359:	ff_dbi <= 8'h40;
		14'h035a:	ff_dbi <= 8'h48;
		14'h035b:	ff_dbi <= 8'h50;
		14'h035c:	ff_dbi <= 8'h60;
		14'h035d:	ff_dbi <= 8'h50;
		14'h035e:	ff_dbi <= 8'h48;
		14'h035f:	ff_dbi <= 8'h00;
		14'h0360:	ff_dbi <= 8'h60;
		14'h0361:	ff_dbi <= 8'h20;
		14'h0362:	ff_dbi <= 8'h20;
		14'h0363:	ff_dbi <= 8'h20;
		14'h0364:	ff_dbi <= 8'h20;
		14'h0365:	ff_dbi <= 8'h20;
		14'h0366:	ff_dbi <= 8'h70;
		14'h0367:	ff_dbi <= 8'h00;
		14'h0368:	ff_dbi <= 8'h00;
		14'h0369:	ff_dbi <= 8'h00;
		14'h036a:	ff_dbi <= 8'hd0;
		14'h036b:	ff_dbi <= 8'ha8;
		14'h036c:	ff_dbi <= 8'ha8;
		14'h036d:	ff_dbi <= 8'ha8;
		14'h036e:	ff_dbi <= 8'ha8;
		14'h036f:	ff_dbi <= 8'h00;
		14'h0370:	ff_dbi <= 8'h00;
		14'h0371:	ff_dbi <= 8'h00;
		14'h0372:	ff_dbi <= 8'hb0;
		14'h0373:	ff_dbi <= 8'hc8;
		14'h0374:	ff_dbi <= 8'h88;
		14'h0375:	ff_dbi <= 8'h88;
		14'h0376:	ff_dbi <= 8'h88;
		14'h0377:	ff_dbi <= 8'h00;
		14'h0378:	ff_dbi <= 8'h00;
		14'h0379:	ff_dbi <= 8'h00;
		14'h037a:	ff_dbi <= 8'h70;
		14'h037b:	ff_dbi <= 8'h88;
		14'h037c:	ff_dbi <= 8'h88;
		14'h037d:	ff_dbi <= 8'h88;
		14'h037e:	ff_dbi <= 8'h70;
		14'h037f:	ff_dbi <= 8'h00;
		14'h0380:	ff_dbi <= 8'h00;
		14'h0381:	ff_dbi <= 8'h00;
		14'h0382:	ff_dbi <= 8'hb0;
		14'h0383:	ff_dbi <= 8'hc8;
		14'h0384:	ff_dbi <= 8'hc8;
		14'h0385:	ff_dbi <= 8'hb0;
		14'h0386:	ff_dbi <= 8'h80;
		14'h0387:	ff_dbi <= 8'h80;
		14'h0388:	ff_dbi <= 8'h00;
		14'h0389:	ff_dbi <= 8'h00;
		14'h038a:	ff_dbi <= 8'h68;
		14'h038b:	ff_dbi <= 8'h98;
		14'h038c:	ff_dbi <= 8'h98;
		14'h038d:	ff_dbi <= 8'h68;
		14'h038e:	ff_dbi <= 8'h08;
		14'h038f:	ff_dbi <= 8'h08;
		14'h0390:	ff_dbi <= 8'h00;
		14'h0391:	ff_dbi <= 8'h00;
		14'h0392:	ff_dbi <= 8'hb0;
		14'h0393:	ff_dbi <= 8'hc8;
		14'h0394:	ff_dbi <= 8'h80;
		14'h0395:	ff_dbi <= 8'h80;
		14'h0396:	ff_dbi <= 8'h80;
		14'h0397:	ff_dbi <= 8'h00;
		14'h0398:	ff_dbi <= 8'h00;
		14'h0399:	ff_dbi <= 8'h00;
		14'h039a:	ff_dbi <= 8'h78;
		14'h039b:	ff_dbi <= 8'h80;
		14'h039c:	ff_dbi <= 8'hf0;
		14'h039d:	ff_dbi <= 8'h08;
		14'h039e:	ff_dbi <= 8'hf0;
		14'h039f:	ff_dbi <= 8'h00;
		14'h03a0:	ff_dbi <= 8'h40;
		14'h03a1:	ff_dbi <= 8'h40;
		14'h03a2:	ff_dbi <= 8'hf0;
		14'h03a3:	ff_dbi <= 8'h40;
		14'h03a4:	ff_dbi <= 8'h40;
		14'h03a5:	ff_dbi <= 8'h48;
		14'h03a6:	ff_dbi <= 8'h30;
		14'h03a7:	ff_dbi <= 8'h00;
		14'h03a8:	ff_dbi <= 8'h00;
		14'h03a9:	ff_dbi <= 8'h00;
		14'h03aa:	ff_dbi <= 8'h90;
		14'h03ab:	ff_dbi <= 8'h90;
		14'h03ac:	ff_dbi <= 8'h90;
		14'h03ad:	ff_dbi <= 8'h90;
		14'h03ae:	ff_dbi <= 8'h68;
		14'h03af:	ff_dbi <= 8'h00;
		14'h03b0:	ff_dbi <= 8'h00;
		14'h03b1:	ff_dbi <= 8'h00;
		14'h03b2:	ff_dbi <= 8'h88;
		14'h03b3:	ff_dbi <= 8'h88;
		14'h03b4:	ff_dbi <= 8'h88;
		14'h03b5:	ff_dbi <= 8'h50;
		14'h03b6:	ff_dbi <= 8'h20;
		14'h03b7:	ff_dbi <= 8'h00;
		14'h03b8:	ff_dbi <= 8'h00;
		14'h03b9:	ff_dbi <= 8'h00;
		14'h03ba:	ff_dbi <= 8'h88;
		14'h03bb:	ff_dbi <= 8'ha8;
		14'h03bc:	ff_dbi <= 8'ha8;
		14'h03bd:	ff_dbi <= 8'ha8;
		14'h03be:	ff_dbi <= 8'h50;
		14'h03bf:	ff_dbi <= 8'h00;
		14'h03c0:	ff_dbi <= 8'h00;
		14'h03c1:	ff_dbi <= 8'h00;
		14'h03c2:	ff_dbi <= 8'h88;
		14'h03c3:	ff_dbi <= 8'h50;
		14'h03c4:	ff_dbi <= 8'h20;
		14'h03c5:	ff_dbi <= 8'h50;
		14'h03c6:	ff_dbi <= 8'h88;
		14'h03c7:	ff_dbi <= 8'h00;
		14'h03c8:	ff_dbi <= 8'h00;
		14'h03c9:	ff_dbi <= 8'h00;
		14'h03ca:	ff_dbi <= 8'h88;
		14'h03cb:	ff_dbi <= 8'h88;
		14'h03cc:	ff_dbi <= 8'h98;
		14'h03cd:	ff_dbi <= 8'h68;
		14'h03ce:	ff_dbi <= 8'h08;
		14'h03cf:	ff_dbi <= 8'h70;
		14'h03d0:	ff_dbi <= 8'h00;
		14'h03d1:	ff_dbi <= 8'h00;
		14'h03d2:	ff_dbi <= 8'hf8;
		14'h03d3:	ff_dbi <= 8'h10;
		14'h03d4:	ff_dbi <= 8'h20;
		14'h03d5:	ff_dbi <= 8'h40;
		14'h03d6:	ff_dbi <= 8'hf8;
		14'h03d7:	ff_dbi <= 8'h00;
		14'h03d8:	ff_dbi <= 8'h18;
		14'h03d9:	ff_dbi <= 8'h20;
		14'h03da:	ff_dbi <= 8'h20;
		14'h03db:	ff_dbi <= 8'h40;
		14'h03dc:	ff_dbi <= 8'h20;
		14'h03dd:	ff_dbi <= 8'h20;
		14'h03de:	ff_dbi <= 8'h18;
		14'h03df:	ff_dbi <= 8'h00;
		14'h03e0:	ff_dbi <= 8'h20;
		14'h03e1:	ff_dbi <= 8'h20;
		14'h03e2:	ff_dbi <= 8'h20;
		14'h03e3:	ff_dbi <= 8'h00;
		14'h03e4:	ff_dbi <= 8'h20;
		14'h03e5:	ff_dbi <= 8'h20;
		14'h03e6:	ff_dbi <= 8'h20;
		14'h03e7:	ff_dbi <= 8'h00;
		14'h03e8:	ff_dbi <= 8'hc0;
		14'h03e9:	ff_dbi <= 8'h20;
		14'h03ea:	ff_dbi <= 8'h20;
		14'h03eb:	ff_dbi <= 8'h10;
		14'h03ec:	ff_dbi <= 8'h20;
		14'h03ed:	ff_dbi <= 8'h20;
		14'h03ee:	ff_dbi <= 8'hc0;
		14'h03ef:	ff_dbi <= 8'h00;
		14'h03f0:	ff_dbi <= 8'h40;
		14'h03f1:	ff_dbi <= 8'ha8;
		14'h03f2:	ff_dbi <= 8'h10;
		14'h03f3:	ff_dbi <= 8'h00;
		14'h03f4:	ff_dbi <= 8'h00;
		14'h03f5:	ff_dbi <= 8'h00;
		14'h03f6:	ff_dbi <= 8'h00;
		14'h03f7:	ff_dbi <= 8'h00;
		14'h03f8:	ff_dbi <= 8'h00;
		14'h03f9:	ff_dbi <= 8'h00;
		14'h03fa:	ff_dbi <= 8'h00;
		14'h03fb:	ff_dbi <= 8'h00;
		14'h03fc:	ff_dbi <= 8'h00;
		14'h03fd:	ff_dbi <= 8'h00;
		14'h03fe:	ff_dbi <= 8'h00;
		14'h03ff:	ff_dbi <= 8'h00;
		14'h0400:	ff_dbi <= 8'h10;
		14'h0401:	ff_dbi <= 8'h38;
		14'h0402:	ff_dbi <= 8'h7c;
		14'h0403:	ff_dbi <= 8'hfe;
		14'h0404:	ff_dbi <= 8'hfe;
		14'h0405:	ff_dbi <= 8'h38;
		14'h0406:	ff_dbi <= 8'h7c;
		14'h0407:	ff_dbi <= 8'h00;
		14'h0408:	ff_dbi <= 8'h6c;
		14'h0409:	ff_dbi <= 8'hfe;
		14'h040a:	ff_dbi <= 8'hfe;
		14'h040b:	ff_dbi <= 8'hfe;
		14'h040c:	ff_dbi <= 8'h7c;
		14'h040d:	ff_dbi <= 8'h38;
		14'h040e:	ff_dbi <= 8'h10;
		14'h040f:	ff_dbi <= 8'h00;
		14'h0410:	ff_dbi <= 8'h38;
		14'h0411:	ff_dbi <= 8'h38;
		14'h0412:	ff_dbi <= 8'hfe;
		14'h0413:	ff_dbi <= 8'hfe;
		14'h0414:	ff_dbi <= 8'hd6;
		14'h0415:	ff_dbi <= 8'h10;
		14'h0416:	ff_dbi <= 8'h7c;
		14'h0417:	ff_dbi <= 8'h00;
		14'h0418:	ff_dbi <= 8'h10;
		14'h0419:	ff_dbi <= 8'h38;
		14'h041a:	ff_dbi <= 8'h7c;
		14'h041b:	ff_dbi <= 8'hfe;
		14'h041c:	ff_dbi <= 8'h7c;
		14'h041d:	ff_dbi <= 8'h38;
		14'h041e:	ff_dbi <= 8'h10;
		14'h041f:	ff_dbi <= 8'h00;
		14'h0420:	ff_dbi <= 8'h00;
		14'h0421:	ff_dbi <= 8'h78;
		14'h0422:	ff_dbi <= 8'h84;
		14'h0423:	ff_dbi <= 8'h84;
		14'h0424:	ff_dbi <= 8'h84;
		14'h0425:	ff_dbi <= 8'h84;
		14'h0426:	ff_dbi <= 8'h78;
		14'h0427:	ff_dbi <= 8'h00;
		14'h0428:	ff_dbi <= 8'h00;
		14'h0429:	ff_dbi <= 8'h78;
		14'h042a:	ff_dbi <= 8'hfc;
		14'h042b:	ff_dbi <= 8'hfc;
		14'h042c:	ff_dbi <= 8'hfc;
		14'h042d:	ff_dbi <= 8'hfc;
		14'h042e:	ff_dbi <= 8'h78;
		14'h042f:	ff_dbi <= 8'h00;
		14'h0430:	ff_dbi <= 8'h20;
		14'h0431:	ff_dbi <= 8'hf0;
		14'h0432:	ff_dbi <= 8'h4c;
		14'h0433:	ff_dbi <= 8'h70;
		14'h0434:	ff_dbi <= 8'ha8;
		14'h0435:	ff_dbi <= 8'h40;
		14'h0436:	ff_dbi <= 8'h3c;
		14'h0437:	ff_dbi <= 8'h00;
		14'h0438:	ff_dbi <= 8'h00;
		14'h0439:	ff_dbi <= 8'h20;
		14'h043a:	ff_dbi <= 8'h78;
		14'h043b:	ff_dbi <= 8'h20;
		14'h043c:	ff_dbi <= 8'h78;
		14'h043d:	ff_dbi <= 8'hb4;
		14'h043e:	ff_dbi <= 8'h64;
		14'h043f:	ff_dbi <= 8'h00;
		14'h0440:	ff_dbi <= 8'h00;
		14'h0441:	ff_dbi <= 8'h00;
		14'h0442:	ff_dbi <= 8'h88;
		14'h0443:	ff_dbi <= 8'h84;
		14'h0444:	ff_dbi <= 8'h84;
		14'h0445:	ff_dbi <= 8'h84;
		14'h0446:	ff_dbi <= 8'h40;
		14'h0447:	ff_dbi <= 8'h00;
		14'h0448:	ff_dbi <= 8'h00;
		14'h0449:	ff_dbi <= 8'h70;
		14'h044a:	ff_dbi <= 8'h00;
		14'h044b:	ff_dbi <= 8'h70;
		14'h044c:	ff_dbi <= 8'h88;
		14'h044d:	ff_dbi <= 8'h08;
		14'h044e:	ff_dbi <= 8'h30;
		14'h044f:	ff_dbi <= 8'h00;
		14'h0450:	ff_dbi <= 8'h00;
		14'h0451:	ff_dbi <= 8'h70;
		14'h0452:	ff_dbi <= 8'h00;
		14'h0453:	ff_dbi <= 8'hf0;
		14'h0454:	ff_dbi <= 8'h20;
		14'h0455:	ff_dbi <= 8'h60;
		14'h0456:	ff_dbi <= 8'h98;
		14'h0457:	ff_dbi <= 8'h00;
		14'h0458:	ff_dbi <= 8'h00;
		14'h0459:	ff_dbi <= 8'h20;
		14'h045a:	ff_dbi <= 8'hf8;
		14'h045b:	ff_dbi <= 8'h24;
		14'h045c:	ff_dbi <= 8'h78;
		14'h045d:	ff_dbi <= 8'ha4;
		14'h045e:	ff_dbi <= 8'h68;
		14'h045f:	ff_dbi <= 8'h00;
		14'h0460:	ff_dbi <= 8'h00;
		14'h0461:	ff_dbi <= 8'h90;
		14'h0462:	ff_dbi <= 8'h58;
		14'h0463:	ff_dbi <= 8'h64;
		14'h0464:	ff_dbi <= 8'ha8;
		14'h0465:	ff_dbi <= 8'h20;
		14'h0466:	ff_dbi <= 8'h10;
		14'h0467:	ff_dbi <= 8'h00;
		14'h0468:	ff_dbi <= 8'h00;
		14'h0469:	ff_dbi <= 8'h10;
		14'h046a:	ff_dbi <= 8'hb8;
		14'h046b:	ff_dbi <= 8'hd4;
		14'h046c:	ff_dbi <= 8'h94;
		14'h046d:	ff_dbi <= 8'h18;
		14'h046e:	ff_dbi <= 8'h20;
		14'h046f:	ff_dbi <= 8'h00;
		14'h0470:	ff_dbi <= 8'h00;
		14'h0471:	ff_dbi <= 8'h10;
		14'h0472:	ff_dbi <= 8'h1c;
		14'h0473:	ff_dbi <= 8'h10;
		14'h0474:	ff_dbi <= 8'h70;
		14'h0475:	ff_dbi <= 8'h98;
		14'h0476:	ff_dbi <= 8'h74;
		14'h0477:	ff_dbi <= 8'h00;
		14'h0478:	ff_dbi <= 8'h00;
		14'h0479:	ff_dbi <= 8'h00;
		14'h047a:	ff_dbi <= 8'h00;
		14'h047b:	ff_dbi <= 8'h78;
		14'h047c:	ff_dbi <= 8'h04;
		14'h047d:	ff_dbi <= 8'h04;
		14'h047e:	ff_dbi <= 8'h38;
		14'h047f:	ff_dbi <= 8'h00;
		14'h0480:	ff_dbi <= 8'h00;
		14'h0481:	ff_dbi <= 8'h00;
		14'h0482:	ff_dbi <= 8'h00;
		14'h0483:	ff_dbi <= 8'h00;
		14'h0484:	ff_dbi <= 8'h00;
		14'h0485:	ff_dbi <= 8'h00;
		14'h0486:	ff_dbi <= 8'h00;
		14'h0487:	ff_dbi <= 8'h00;
		14'h0488:	ff_dbi <= 8'h20;
		14'h0489:	ff_dbi <= 8'h7c;
		14'h048a:	ff_dbi <= 8'h20;
		14'h048b:	ff_dbi <= 8'h7c;
		14'h048c:	ff_dbi <= 8'haa;
		14'h048d:	ff_dbi <= 8'h92;
		14'h048e:	ff_dbi <= 8'h64;
		14'h048f:	ff_dbi <= 8'h00;
		14'h0490:	ff_dbi <= 8'h00;
		14'h0491:	ff_dbi <= 8'h84;
		14'h0492:	ff_dbi <= 8'h82;
		14'h0493:	ff_dbi <= 8'h82;
		14'h0494:	ff_dbi <= 8'h82;
		14'h0495:	ff_dbi <= 8'h80;
		14'h0496:	ff_dbi <= 8'h40;
		14'h0497:	ff_dbi <= 8'h00;
		14'h0498:	ff_dbi <= 8'h38;
		14'h0499:	ff_dbi <= 8'h00;
		14'h049a:	ff_dbi <= 8'h38;
		14'h049b:	ff_dbi <= 8'h44;
		14'h049c:	ff_dbi <= 8'h04;
		14'h049d:	ff_dbi <= 8'h08;
		14'h049e:	ff_dbi <= 8'h30;
		14'h049f:	ff_dbi <= 8'h00;
		14'h04a0:	ff_dbi <= 8'h70;
		14'h04a1:	ff_dbi <= 8'h00;
		14'h04a2:	ff_dbi <= 8'hf8;
		14'h04a3:	ff_dbi <= 8'h10;
		14'h04a4:	ff_dbi <= 8'h20;
		14'h04a5:	ff_dbi <= 8'h60;
		14'h04a6:	ff_dbi <= 8'h9c;
		14'h04a7:	ff_dbi <= 8'h00;
		14'h04a8:	ff_dbi <= 8'h24;
		14'h04a9:	ff_dbi <= 8'hfa;
		14'h04aa:	ff_dbi <= 8'h20;
		14'h04ab:	ff_dbi <= 8'h7c;
		14'h04ac:	ff_dbi <= 8'ha2;
		14'h04ad:	ff_dbi <= 8'ha2;
		14'h04ae:	ff_dbi <= 8'h44;
		14'h04af:	ff_dbi <= 8'h00;
		14'h04b0:	ff_dbi <= 8'h40;
		14'h04b1:	ff_dbi <= 8'h44;
		14'h04b2:	ff_dbi <= 8'hf2;
		14'h04b3:	ff_dbi <= 8'h4a;
		14'h04b4:	ff_dbi <= 8'h48;
		14'h04b5:	ff_dbi <= 8'h88;
		14'h04b6:	ff_dbi <= 8'h30;
		14'h04b7:	ff_dbi <= 8'h00;
		14'h04b8:	ff_dbi <= 8'h20;
		14'h04b9:	ff_dbi <= 8'hfc;
		14'h04ba:	ff_dbi <= 8'h10;
		14'h04bb:	ff_dbi <= 8'hfc;
		14'h04bc:	ff_dbi <= 8'h08;
		14'h04bd:	ff_dbi <= 8'h80;
		14'h04be:	ff_dbi <= 8'h78;
		14'h04bf:	ff_dbi <= 8'h00;
		14'h04c0:	ff_dbi <= 8'h08;
		14'h04c1:	ff_dbi <= 8'h10;
		14'h04c2:	ff_dbi <= 8'h20;
		14'h04c3:	ff_dbi <= 8'h40;
		14'h04c4:	ff_dbi <= 8'h20;
		14'h04c5:	ff_dbi <= 8'h10;
		14'h04c6:	ff_dbi <= 8'h08;
		14'h04c7:	ff_dbi <= 8'h00;
		14'h04c8:	ff_dbi <= 8'h04;
		14'h04c9:	ff_dbi <= 8'h84;
		14'h04ca:	ff_dbi <= 8'h9e;
		14'h04cb:	ff_dbi <= 8'h84;
		14'h04cc:	ff_dbi <= 8'h84;
		14'h04cd:	ff_dbi <= 8'h84;
		14'h04ce:	ff_dbi <= 8'h48;
		14'h04cf:	ff_dbi <= 8'h00;
		14'h04d0:	ff_dbi <= 8'h78;
		14'h04d1:	ff_dbi <= 8'h04;
		14'h04d2:	ff_dbi <= 8'h00;
		14'h04d3:	ff_dbi <= 8'h00;
		14'h04d4:	ff_dbi <= 8'h00;
		14'h04d5:	ff_dbi <= 8'h80;
		14'h04d6:	ff_dbi <= 8'h7c;
		14'h04d7:	ff_dbi <= 8'h00;
		14'h04d8:	ff_dbi <= 8'h10;
		14'h04d9:	ff_dbi <= 8'hfe;
		14'h04da:	ff_dbi <= 8'h08;
		14'h04db:	ff_dbi <= 8'h04;
		14'h04dc:	ff_dbi <= 8'h04;
		14'h04dd:	ff_dbi <= 8'h80;
		14'h04de:	ff_dbi <= 8'h78;
		14'h04df:	ff_dbi <= 8'h00;
		14'h04e0:	ff_dbi <= 8'h80;
		14'h04e1:	ff_dbi <= 8'h80;
		14'h04e2:	ff_dbi <= 8'h80;
		14'h04e3:	ff_dbi <= 8'h80;
		14'h04e4:	ff_dbi <= 8'h84;
		14'h04e5:	ff_dbi <= 8'h88;
		14'h04e6:	ff_dbi <= 8'h70;
		14'h04e7:	ff_dbi <= 8'h00;
		14'h04e8:	ff_dbi <= 8'h08;
		14'h04e9:	ff_dbi <= 8'hfe;
		14'h04ea:	ff_dbi <= 8'h38;
		14'h04eb:	ff_dbi <= 8'h48;
		14'h04ec:	ff_dbi <= 8'h38;
		14'h04ed:	ff_dbi <= 8'h08;
		14'h04ee:	ff_dbi <= 8'h10;
		14'h04ef:	ff_dbi <= 8'h00;
		14'h04f0:	ff_dbi <= 8'h44;
		14'h04f1:	ff_dbi <= 8'h44;
		14'h04f2:	ff_dbi <= 8'hfe;
		14'h04f3:	ff_dbi <= 8'h44;
		14'h04f4:	ff_dbi <= 8'h48;
		14'h04f5:	ff_dbi <= 8'h40;
		14'h04f6:	ff_dbi <= 8'h3c;
		14'h04f7:	ff_dbi <= 8'h00;
		14'h04f8:	ff_dbi <= 8'h44;
		14'h04f9:	ff_dbi <= 8'h28;
		14'h04fa:	ff_dbi <= 8'hfe;
		14'h04fb:	ff_dbi <= 8'h20;
		14'h04fc:	ff_dbi <= 8'h40;
		14'h04fd:	ff_dbi <= 8'h40;
		14'h04fe:	ff_dbi <= 8'h3c;
		14'h04ff:	ff_dbi <= 8'h00;
		14'h0500:	ff_dbi <= 8'h00;
		14'h0501:	ff_dbi <= 8'h00;
		14'h0502:	ff_dbi <= 8'h00;
		14'h0503:	ff_dbi <= 8'h00;
		14'h0504:	ff_dbi <= 8'h00;
		14'h0505:	ff_dbi <= 8'h00;
		14'h0506:	ff_dbi <= 8'h00;
		14'h0507:	ff_dbi <= 8'h00;
		14'h0508:	ff_dbi <= 8'h00;
		14'h0509:	ff_dbi <= 8'h00;
		14'h050a:	ff_dbi <= 8'h00;
		14'h050b:	ff_dbi <= 8'h00;
		14'h050c:	ff_dbi <= 8'h60;
		14'h050d:	ff_dbi <= 8'h90;
		14'h050e:	ff_dbi <= 8'h60;
		14'h050f:	ff_dbi <= 8'h00;
		14'h0510:	ff_dbi <= 8'h38;
		14'h0511:	ff_dbi <= 8'h20;
		14'h0512:	ff_dbi <= 8'h20;
		14'h0513:	ff_dbi <= 8'h20;
		14'h0514:	ff_dbi <= 8'h00;
		14'h0515:	ff_dbi <= 8'h00;
		14'h0516:	ff_dbi <= 8'h00;
		14'h0517:	ff_dbi <= 8'h00;
		14'h0518:	ff_dbi <= 8'h00;
		14'h0519:	ff_dbi <= 8'h00;
		14'h051a:	ff_dbi <= 8'h00;
		14'h051b:	ff_dbi <= 8'h20;
		14'h051c:	ff_dbi <= 8'h20;
		14'h051d:	ff_dbi <= 8'h20;
		14'h051e:	ff_dbi <= 8'he0;
		14'h051f:	ff_dbi <= 8'h00;
		14'h0520:	ff_dbi <= 8'h00;
		14'h0521:	ff_dbi <= 8'h00;
		14'h0522:	ff_dbi <= 8'h00;
		14'h0523:	ff_dbi <= 8'h00;
		14'h0524:	ff_dbi <= 8'h80;
		14'h0525:	ff_dbi <= 8'h40;
		14'h0526:	ff_dbi <= 8'h20;
		14'h0527:	ff_dbi <= 8'h00;
		14'h0528:	ff_dbi <= 8'h00;
		14'h0529:	ff_dbi <= 8'h00;
		14'h052a:	ff_dbi <= 8'h00;
		14'h052b:	ff_dbi <= 8'h30;
		14'h052c:	ff_dbi <= 8'h30;
		14'h052d:	ff_dbi <= 8'h00;
		14'h052e:	ff_dbi <= 8'h00;
		14'h052f:	ff_dbi <= 8'h00;
		14'h0530:	ff_dbi <= 8'hf8;
		14'h0531:	ff_dbi <= 8'h08;
		14'h0532:	ff_dbi <= 8'hf8;
		14'h0533:	ff_dbi <= 8'h08;
		14'h0534:	ff_dbi <= 8'h10;
		14'h0535:	ff_dbi <= 8'h20;
		14'h0536:	ff_dbi <= 8'h40;
		14'h0537:	ff_dbi <= 8'h00;
		14'h0538:	ff_dbi <= 8'h00;
		14'h0539:	ff_dbi <= 8'h00;
		14'h053a:	ff_dbi <= 8'hf0;
		14'h053b:	ff_dbi <= 8'h10;
		14'h053c:	ff_dbi <= 8'h60;
		14'h053d:	ff_dbi <= 8'h40;
		14'h053e:	ff_dbi <= 8'h80;
		14'h053f:	ff_dbi <= 8'h00;
		14'h0540:	ff_dbi <= 8'h00;
		14'h0541:	ff_dbi <= 8'h10;
		14'h0542:	ff_dbi <= 8'h20;
		14'h0543:	ff_dbi <= 8'h60;
		14'h0544:	ff_dbi <= 8'ha0;
		14'h0545:	ff_dbi <= 8'h20;
		14'h0546:	ff_dbi <= 8'h20;
		14'h0547:	ff_dbi <= 8'h00;
		14'h0548:	ff_dbi <= 8'h00;
		14'h0549:	ff_dbi <= 8'h20;
		14'h054a:	ff_dbi <= 8'hf0;
		14'h054b:	ff_dbi <= 8'h90;
		14'h054c:	ff_dbi <= 8'h10;
		14'h054d:	ff_dbi <= 8'h20;
		14'h054e:	ff_dbi <= 8'h40;
		14'h054f:	ff_dbi <= 8'h00;
		14'h0550:	ff_dbi <= 8'h00;
		14'h0551:	ff_dbi <= 8'h00;
		14'h0552:	ff_dbi <= 8'hf0;
		14'h0553:	ff_dbi <= 8'h20;
		14'h0554:	ff_dbi <= 8'h20;
		14'h0555:	ff_dbi <= 8'h20;
		14'h0556:	ff_dbi <= 8'hf0;
		14'h0557:	ff_dbi <= 8'h00;
		14'h0558:	ff_dbi <= 8'h00;
		14'h0559:	ff_dbi <= 8'h20;
		14'h055a:	ff_dbi <= 8'hf0;
		14'h055b:	ff_dbi <= 8'h60;
		14'h055c:	ff_dbi <= 8'ha0;
		14'h055d:	ff_dbi <= 8'ha0;
		14'h055e:	ff_dbi <= 8'h20;
		14'h055f:	ff_dbi <= 8'h00;
		14'h0560:	ff_dbi <= 8'h00;
		14'h0561:	ff_dbi <= 8'h40;
		14'h0562:	ff_dbi <= 8'hf8;
		14'h0563:	ff_dbi <= 8'h48;
		14'h0564:	ff_dbi <= 8'h50;
		14'h0565:	ff_dbi <= 8'h40;
		14'h0566:	ff_dbi <= 8'h40;
		14'h0567:	ff_dbi <= 8'h00;
		14'h0568:	ff_dbi <= 8'h00;
		14'h0569:	ff_dbi <= 8'h00;
		14'h056a:	ff_dbi <= 8'h70;
		14'h056b:	ff_dbi <= 8'h10;
		14'h056c:	ff_dbi <= 8'h10;
		14'h056d:	ff_dbi <= 8'h10;
		14'h056e:	ff_dbi <= 8'hf8;
		14'h056f:	ff_dbi <= 8'h00;
		14'h0570:	ff_dbi <= 8'h00;
		14'h0571:	ff_dbi <= 8'h00;
		14'h0572:	ff_dbi <= 8'hf0;
		14'h0573:	ff_dbi <= 8'h10;
		14'h0574:	ff_dbi <= 8'hf0;
		14'h0575:	ff_dbi <= 8'h10;
		14'h0576:	ff_dbi <= 8'hf0;
		14'h0577:	ff_dbi <= 8'h00;
		14'h0578:	ff_dbi <= 8'h00;
		14'h0579:	ff_dbi <= 8'h00;
		14'h057a:	ff_dbi <= 8'ha8;
		14'h057b:	ff_dbi <= 8'ha8;
		14'h057c:	ff_dbi <= 8'h08;
		14'h057d:	ff_dbi <= 8'h10;
		14'h057e:	ff_dbi <= 8'h20;
		14'h057f:	ff_dbi <= 8'h00;
		14'h0580:	ff_dbi <= 8'h00;
		14'h0581:	ff_dbi <= 8'h00;
		14'h0582:	ff_dbi <= 8'h80;
		14'h0583:	ff_dbi <= 8'h7c;
		14'h0584:	ff_dbi <= 8'h00;
		14'h0585:	ff_dbi <= 8'h00;
		14'h0586:	ff_dbi <= 8'h00;
		14'h0587:	ff_dbi <= 8'h00;
		14'h0588:	ff_dbi <= 8'hf8;
		14'h0589:	ff_dbi <= 8'h08;
		14'h058a:	ff_dbi <= 8'h28;
		14'h058b:	ff_dbi <= 8'h30;
		14'h058c:	ff_dbi <= 8'h20;
		14'h058d:	ff_dbi <= 8'h20;
		14'h058e:	ff_dbi <= 8'h40;
		14'h058f:	ff_dbi <= 8'h00;
		14'h0590:	ff_dbi <= 8'h08;
		14'h0591:	ff_dbi <= 8'h10;
		14'h0592:	ff_dbi <= 8'h20;
		14'h0593:	ff_dbi <= 8'h60;
		14'h0594:	ff_dbi <= 8'ha0;
		14'h0595:	ff_dbi <= 8'h20;
		14'h0596:	ff_dbi <= 8'h20;
		14'h0597:	ff_dbi <= 8'h00;
		14'h0598:	ff_dbi <= 8'h20;
		14'h0599:	ff_dbi <= 8'hf8;
		14'h059a:	ff_dbi <= 8'h88;
		14'h059b:	ff_dbi <= 8'h88;
		14'h059c:	ff_dbi <= 8'h08;
		14'h059d:	ff_dbi <= 8'h10;
		14'h059e:	ff_dbi <= 8'h20;
		14'h059f:	ff_dbi <= 8'h00;
		14'h05a0:	ff_dbi <= 8'h00;
		14'h05a1:	ff_dbi <= 8'hf8;
		14'h05a2:	ff_dbi <= 8'h20;
		14'h05a3:	ff_dbi <= 8'h20;
		14'h05a4:	ff_dbi <= 8'h20;
		14'h05a5:	ff_dbi <= 8'h20;
		14'h05a6:	ff_dbi <= 8'hf8;
		14'h05a7:	ff_dbi <= 8'h00;
		14'h05a8:	ff_dbi <= 8'h10;
		14'h05a9:	ff_dbi <= 8'hf8;
		14'h05aa:	ff_dbi <= 8'h10;
		14'h05ab:	ff_dbi <= 8'h30;
		14'h05ac:	ff_dbi <= 8'h50;
		14'h05ad:	ff_dbi <= 8'h90;
		14'h05ae:	ff_dbi <= 8'h10;
		14'h05af:	ff_dbi <= 8'h00;
		14'h05b0:	ff_dbi <= 8'h20;
		14'h05b1:	ff_dbi <= 8'hf8;
		14'h05b2:	ff_dbi <= 8'h28;
		14'h05b3:	ff_dbi <= 8'h28;
		14'h05b4:	ff_dbi <= 8'h28;
		14'h05b5:	ff_dbi <= 8'h48;
		14'h05b6:	ff_dbi <= 8'h88;
		14'h05b7:	ff_dbi <= 8'h00;
		14'h05b8:	ff_dbi <= 8'h20;
		14'h05b9:	ff_dbi <= 8'hf8;
		14'h05ba:	ff_dbi <= 8'h20;
		14'h05bb:	ff_dbi <= 8'hf8;
		14'h05bc:	ff_dbi <= 8'h20;
		14'h05bd:	ff_dbi <= 8'h20;
		14'h05be:	ff_dbi <= 8'h20;
		14'h05bf:	ff_dbi <= 8'h00;
		14'h05c0:	ff_dbi <= 8'h78;
		14'h05c1:	ff_dbi <= 8'h48;
		14'h05c2:	ff_dbi <= 8'h88;
		14'h05c3:	ff_dbi <= 8'h08;
		14'h05c4:	ff_dbi <= 8'h08;
		14'h05c5:	ff_dbi <= 8'h10;
		14'h05c6:	ff_dbi <= 8'h20;
		14'h05c7:	ff_dbi <= 8'h00;
		14'h05c8:	ff_dbi <= 8'h40;
		14'h05c9:	ff_dbi <= 8'h78;
		14'h05ca:	ff_dbi <= 8'h50;
		14'h05cb:	ff_dbi <= 8'h90;
		14'h05cc:	ff_dbi <= 8'h10;
		14'h05cd:	ff_dbi <= 8'h10;
		14'h05ce:	ff_dbi <= 8'h20;
		14'h05cf:	ff_dbi <= 8'h00;
		14'h05d0:	ff_dbi <= 8'h00;
		14'h05d1:	ff_dbi <= 8'hf8;
		14'h05d2:	ff_dbi <= 8'h08;
		14'h05d3:	ff_dbi <= 8'h08;
		14'h05d4:	ff_dbi <= 8'h08;
		14'h05d5:	ff_dbi <= 8'h08;
		14'h05d6:	ff_dbi <= 8'hf8;
		14'h05d7:	ff_dbi <= 8'h00;
		14'h05d8:	ff_dbi <= 8'h50;
		14'h05d9:	ff_dbi <= 8'hf8;
		14'h05da:	ff_dbi <= 8'h50;
		14'h05db:	ff_dbi <= 8'h50;
		14'h05dc:	ff_dbi <= 8'h10;
		14'h05dd:	ff_dbi <= 8'h10;
		14'h05de:	ff_dbi <= 8'h20;
		14'h05df:	ff_dbi <= 8'h00;
		14'h05e0:	ff_dbi <= 8'h00;
		14'h05e1:	ff_dbi <= 8'hc0;
		14'h05e2:	ff_dbi <= 8'h08;
		14'h05e3:	ff_dbi <= 8'hc8;
		14'h05e4:	ff_dbi <= 8'h08;
		14'h05e5:	ff_dbi <= 8'h10;
		14'h05e6:	ff_dbi <= 8'he0;
		14'h05e7:	ff_dbi <= 8'h00;
		14'h05e8:	ff_dbi <= 8'h00;
		14'h05e9:	ff_dbi <= 8'hf8;
		14'h05ea:	ff_dbi <= 8'h08;
		14'h05eb:	ff_dbi <= 8'h10;
		14'h05ec:	ff_dbi <= 8'h20;
		14'h05ed:	ff_dbi <= 8'h50;
		14'h05ee:	ff_dbi <= 8'h88;
		14'h05ef:	ff_dbi <= 8'h00;
		14'h05f0:	ff_dbi <= 8'h40;
		14'h05f1:	ff_dbi <= 8'hf8;
		14'h05f2:	ff_dbi <= 8'h48;
		14'h05f3:	ff_dbi <= 8'h50;
		14'h05f4:	ff_dbi <= 8'h40;
		14'h05f5:	ff_dbi <= 8'h40;
		14'h05f6:	ff_dbi <= 8'h38;
		14'h05f7:	ff_dbi <= 8'h00;
		14'h05f8:	ff_dbi <= 8'h88;
		14'h05f9:	ff_dbi <= 8'h88;
		14'h05fa:	ff_dbi <= 8'h48;
		14'h05fb:	ff_dbi <= 8'h08;
		14'h05fc:	ff_dbi <= 8'h10;
		14'h05fd:	ff_dbi <= 8'h20;
		14'h05fe:	ff_dbi <= 8'h40;
		14'h05ff:	ff_dbi <= 8'h00;
		14'h0600:	ff_dbi <= 8'h78;
		14'h0601:	ff_dbi <= 8'h48;
		14'h0602:	ff_dbi <= 8'h78;
		14'h0603:	ff_dbi <= 8'h88;
		14'h0604:	ff_dbi <= 8'h08;
		14'h0605:	ff_dbi <= 8'h10;
		14'h0606:	ff_dbi <= 8'h20;
		14'h0607:	ff_dbi <= 8'h00;
		14'h0608:	ff_dbi <= 8'h10;
		14'h0609:	ff_dbi <= 8'he0;
		14'h060a:	ff_dbi <= 8'h20;
		14'h060b:	ff_dbi <= 8'hf8;
		14'h060c:	ff_dbi <= 8'h20;
		14'h060d:	ff_dbi <= 8'h20;
		14'h060e:	ff_dbi <= 8'h40;
		14'h060f:	ff_dbi <= 8'h00;
		14'h0610:	ff_dbi <= 8'ha8;
		14'h0611:	ff_dbi <= 8'ha8;
		14'h0612:	ff_dbi <= 8'ha8;
		14'h0613:	ff_dbi <= 8'h08;
		14'h0614:	ff_dbi <= 8'h08;
		14'h0615:	ff_dbi <= 8'h10;
		14'h0616:	ff_dbi <= 8'h20;
		14'h0617:	ff_dbi <= 8'h00;
		14'h0618:	ff_dbi <= 8'h70;
		14'h0619:	ff_dbi <= 8'h00;
		14'h061a:	ff_dbi <= 8'hf8;
		14'h061b:	ff_dbi <= 8'h20;
		14'h061c:	ff_dbi <= 8'h20;
		14'h061d:	ff_dbi <= 8'h20;
		14'h061e:	ff_dbi <= 8'h40;
		14'h061f:	ff_dbi <= 8'h00;
		14'h0620:	ff_dbi <= 8'h40;
		14'h0621:	ff_dbi <= 8'h40;
		14'h0622:	ff_dbi <= 8'h60;
		14'h0623:	ff_dbi <= 8'h50;
		14'h0624:	ff_dbi <= 8'h48;
		14'h0625:	ff_dbi <= 8'h40;
		14'h0626:	ff_dbi <= 8'h40;
		14'h0627:	ff_dbi <= 8'h00;
		14'h0628:	ff_dbi <= 8'h20;
		14'h0629:	ff_dbi <= 8'hf8;
		14'h062a:	ff_dbi <= 8'h20;
		14'h062b:	ff_dbi <= 8'h20;
		14'h062c:	ff_dbi <= 8'h20;
		14'h062d:	ff_dbi <= 8'h20;
		14'h062e:	ff_dbi <= 8'h40;
		14'h062f:	ff_dbi <= 8'h00;
		14'h0630:	ff_dbi <= 8'h00;
		14'h0631:	ff_dbi <= 8'h70;
		14'h0632:	ff_dbi <= 8'h00;
		14'h0633:	ff_dbi <= 8'h00;
		14'h0634:	ff_dbi <= 8'h00;
		14'h0635:	ff_dbi <= 8'h00;
		14'h0636:	ff_dbi <= 8'hf8;
		14'h0637:	ff_dbi <= 8'h00;
		14'h0638:	ff_dbi <= 8'h00;
		14'h0639:	ff_dbi <= 8'hf8;
		14'h063a:	ff_dbi <= 8'h08;
		14'h063b:	ff_dbi <= 8'hd0;
		14'h063c:	ff_dbi <= 8'h20;
		14'h063d:	ff_dbi <= 8'h50;
		14'h063e:	ff_dbi <= 8'h88;
		14'h063f:	ff_dbi <= 8'h00;
		14'h0640:	ff_dbi <= 8'h20;
		14'h0641:	ff_dbi <= 8'hf8;
		14'h0642:	ff_dbi <= 8'h08;
		14'h0643:	ff_dbi <= 8'h30;
		14'h0644:	ff_dbi <= 8'he8;
		14'h0645:	ff_dbi <= 8'h20;
		14'h0646:	ff_dbi <= 8'h20;
		14'h0647:	ff_dbi <= 8'h00;
		14'h0648:	ff_dbi <= 8'h08;
		14'h0649:	ff_dbi <= 8'h08;
		14'h064a:	ff_dbi <= 8'h08;
		14'h064b:	ff_dbi <= 8'h10;
		14'h064c:	ff_dbi <= 8'h20;
		14'h064d:	ff_dbi <= 8'h40;
		14'h064e:	ff_dbi <= 8'h80;
		14'h064f:	ff_dbi <= 8'h00;
		14'h0650:	ff_dbi <= 8'h20;
		14'h0651:	ff_dbi <= 8'h10;
		14'h0652:	ff_dbi <= 8'h48;
		14'h0653:	ff_dbi <= 8'h48;
		14'h0654:	ff_dbi <= 8'h48;
		14'h0655:	ff_dbi <= 8'h48;
		14'h0656:	ff_dbi <= 8'h88;
		14'h0657:	ff_dbi <= 8'h00;
		14'h0658:	ff_dbi <= 8'h80;
		14'h0659:	ff_dbi <= 8'h80;
		14'h065a:	ff_dbi <= 8'hf8;
		14'h065b:	ff_dbi <= 8'h80;
		14'h065c:	ff_dbi <= 8'h80;
		14'h065d:	ff_dbi <= 8'h80;
		14'h065e:	ff_dbi <= 8'h78;
		14'h065f:	ff_dbi <= 8'h00;
		14'h0660:	ff_dbi <= 8'hf8;
		14'h0661:	ff_dbi <= 8'h08;
		14'h0662:	ff_dbi <= 8'h08;
		14'h0663:	ff_dbi <= 8'h08;
		14'h0664:	ff_dbi <= 8'h10;
		14'h0665:	ff_dbi <= 8'h20;
		14'h0666:	ff_dbi <= 8'h40;
		14'h0667:	ff_dbi <= 8'h00;
		14'h0668:	ff_dbi <= 8'h00;
		14'h0669:	ff_dbi <= 8'h40;
		14'h066a:	ff_dbi <= 8'ha0;
		14'h066b:	ff_dbi <= 8'h10;
		14'h066c:	ff_dbi <= 8'h08;
		14'h066d:	ff_dbi <= 8'h08;
		14'h066e:	ff_dbi <= 8'h00;
		14'h066f:	ff_dbi <= 8'h00;
		14'h0670:	ff_dbi <= 8'h20;
		14'h0671:	ff_dbi <= 8'hf8;
		14'h0672:	ff_dbi <= 8'h20;
		14'h0673:	ff_dbi <= 8'h20;
		14'h0674:	ff_dbi <= 8'ha8;
		14'h0675:	ff_dbi <= 8'ha8;
		14'h0676:	ff_dbi <= 8'h20;
		14'h0677:	ff_dbi <= 8'h00;
		14'h0678:	ff_dbi <= 8'h00;
		14'h0679:	ff_dbi <= 8'hf8;
		14'h067a:	ff_dbi <= 8'h08;
		14'h067b:	ff_dbi <= 8'h08;
		14'h067c:	ff_dbi <= 8'h50;
		14'h067d:	ff_dbi <= 8'h20;
		14'h067e:	ff_dbi <= 8'h10;
		14'h067f:	ff_dbi <= 8'h00;
		14'h0680:	ff_dbi <= 8'hf0;
		14'h0681:	ff_dbi <= 8'h00;
		14'h0682:	ff_dbi <= 8'h60;
		14'h0683:	ff_dbi <= 8'h00;
		14'h0684:	ff_dbi <= 8'h00;
		14'h0685:	ff_dbi <= 8'hf0;
		14'h0686:	ff_dbi <= 8'h08;
		14'h0687:	ff_dbi <= 8'h00;
		14'h0688:	ff_dbi <= 8'h10;
		14'h0689:	ff_dbi <= 8'h20;
		14'h068a:	ff_dbi <= 8'h40;
		14'h068b:	ff_dbi <= 8'h80;
		14'h068c:	ff_dbi <= 8'h90;
		14'h068d:	ff_dbi <= 8'h88;
		14'h068e:	ff_dbi <= 8'hf8;
		14'h068f:	ff_dbi <= 8'h00;
		14'h0690:	ff_dbi <= 8'h08;
		14'h0691:	ff_dbi <= 8'h08;
		14'h0692:	ff_dbi <= 8'h08;
		14'h0693:	ff_dbi <= 8'h50;
		14'h0694:	ff_dbi <= 8'h20;
		14'h0695:	ff_dbi <= 8'h50;
		14'h0696:	ff_dbi <= 8'h80;
		14'h0697:	ff_dbi <= 8'h00;
		14'h0698:	ff_dbi <= 8'h78;
		14'h0699:	ff_dbi <= 8'h20;
		14'h069a:	ff_dbi <= 8'hf8;
		14'h069b:	ff_dbi <= 8'h20;
		14'h069c:	ff_dbi <= 8'h20;
		14'h069d:	ff_dbi <= 8'h20;
		14'h069e:	ff_dbi <= 8'h18;
		14'h069f:	ff_dbi <= 8'h00;
		14'h06a0:	ff_dbi <= 8'h40;
		14'h06a1:	ff_dbi <= 8'hf8;
		14'h06a2:	ff_dbi <= 8'h48;
		14'h06a3:	ff_dbi <= 8'h48;
		14'h06a4:	ff_dbi <= 8'h50;
		14'h06a5:	ff_dbi <= 8'h40;
		14'h06a6:	ff_dbi <= 8'h40;
		14'h06a7:	ff_dbi <= 8'h00;
		14'h06a8:	ff_dbi <= 8'h00;
		14'h06a9:	ff_dbi <= 8'h70;
		14'h06aa:	ff_dbi <= 8'h10;
		14'h06ab:	ff_dbi <= 8'h10;
		14'h06ac:	ff_dbi <= 8'h10;
		14'h06ad:	ff_dbi <= 8'h10;
		14'h06ae:	ff_dbi <= 8'hf8;
		14'h06af:	ff_dbi <= 8'h00;
		14'h06b0:	ff_dbi <= 8'h00;
		14'h06b1:	ff_dbi <= 8'hf8;
		14'h06b2:	ff_dbi <= 8'h08;
		14'h06b3:	ff_dbi <= 8'hf8;
		14'h06b4:	ff_dbi <= 8'h08;
		14'h06b5:	ff_dbi <= 8'h08;
		14'h06b6:	ff_dbi <= 8'hf8;
		14'h06b7:	ff_dbi <= 8'h00;
		14'h06b8:	ff_dbi <= 8'h70;
		14'h06b9:	ff_dbi <= 8'h00;
		14'h06ba:	ff_dbi <= 8'hf8;
		14'h06bb:	ff_dbi <= 8'h08;
		14'h06bc:	ff_dbi <= 8'h08;
		14'h06bd:	ff_dbi <= 8'h10;
		14'h06be:	ff_dbi <= 8'h20;
		14'h06bf:	ff_dbi <= 8'h00;
		14'h06c0:	ff_dbi <= 8'h48;
		14'h06c1:	ff_dbi <= 8'h48;
		14'h06c2:	ff_dbi <= 8'h48;
		14'h06c3:	ff_dbi <= 8'h48;
		14'h06c4:	ff_dbi <= 8'h48;
		14'h06c5:	ff_dbi <= 8'h10;
		14'h06c6:	ff_dbi <= 8'h20;
		14'h06c7:	ff_dbi <= 8'h00;
		14'h06c8:	ff_dbi <= 8'h10;
		14'h06c9:	ff_dbi <= 8'h50;
		14'h06ca:	ff_dbi <= 8'h50;
		14'h06cb:	ff_dbi <= 8'h50;
		14'h06cc:	ff_dbi <= 8'h50;
		14'h06cd:	ff_dbi <= 8'h58;
		14'h06ce:	ff_dbi <= 8'h90;
		14'h06cf:	ff_dbi <= 8'h00;
		14'h06d0:	ff_dbi <= 8'h40;
		14'h06d1:	ff_dbi <= 8'h40;
		14'h06d2:	ff_dbi <= 8'h40;
		14'h06d3:	ff_dbi <= 8'h48;
		14'h06d4:	ff_dbi <= 8'h48;
		14'h06d5:	ff_dbi <= 8'h50;
		14'h06d6:	ff_dbi <= 8'h60;
		14'h06d7:	ff_dbi <= 8'h00;
		14'h06d8:	ff_dbi <= 8'h00;
		14'h06d9:	ff_dbi <= 8'hf8;
		14'h06da:	ff_dbi <= 8'h88;
		14'h06db:	ff_dbi <= 8'h88;
		14'h06dc:	ff_dbi <= 8'h88;
		14'h06dd:	ff_dbi <= 8'h88;
		14'h06de:	ff_dbi <= 8'hf8;
		14'h06df:	ff_dbi <= 8'h00;
		14'h06e0:	ff_dbi <= 8'hf8;
		14'h06e1:	ff_dbi <= 8'h88;
		14'h06e2:	ff_dbi <= 8'h88;
		14'h06e3:	ff_dbi <= 8'h08;
		14'h06e4:	ff_dbi <= 8'h08;
		14'h06e5:	ff_dbi <= 8'h10;
		14'h06e6:	ff_dbi <= 8'h20;
		14'h06e7:	ff_dbi <= 8'h00;
		14'h06e8:	ff_dbi <= 8'h00;
		14'h06e9:	ff_dbi <= 8'hc0;
		14'h06ea:	ff_dbi <= 8'h00;
		14'h06eb:	ff_dbi <= 8'h08;
		14'h06ec:	ff_dbi <= 8'h08;
		14'h06ed:	ff_dbi <= 8'h10;
		14'h06ee:	ff_dbi <= 8'he0;
		14'h06ef:	ff_dbi <= 8'h00;
		14'h06f0:	ff_dbi <= 8'h90;
		14'h06f1:	ff_dbi <= 8'h48;
		14'h06f2:	ff_dbi <= 8'h00;
		14'h06f3:	ff_dbi <= 8'h00;
		14'h06f4:	ff_dbi <= 8'h00;
		14'h06f5:	ff_dbi <= 8'h00;
		14'h06f6:	ff_dbi <= 8'h00;
		14'h06f7:	ff_dbi <= 8'h00;
		14'h06f8:	ff_dbi <= 8'h60;
		14'h06f9:	ff_dbi <= 8'h90;
		14'h06fa:	ff_dbi <= 8'h60;
		14'h06fb:	ff_dbi <= 8'h00;
		14'h06fc:	ff_dbi <= 8'h00;
		14'h06fd:	ff_dbi <= 8'h00;
		14'h06fe:	ff_dbi <= 8'h00;
		14'h06ff:	ff_dbi <= 8'h00;
		14'h0700:	ff_dbi <= 8'h20;
		14'h0701:	ff_dbi <= 8'hf8;
		14'h0702:	ff_dbi <= 8'h20;
		14'h0703:	ff_dbi <= 8'h4e;
		14'h0704:	ff_dbi <= 8'h40;
		14'h0705:	ff_dbi <= 8'h90;
		14'h0706:	ff_dbi <= 8'h8e;
		14'h0707:	ff_dbi <= 8'h00;
		14'h0708:	ff_dbi <= 8'h10;
		14'h0709:	ff_dbi <= 8'hfe;
		14'h070a:	ff_dbi <= 8'h20;
		14'h070b:	ff_dbi <= 8'h78;
		14'h070c:	ff_dbi <= 8'h04;
		14'h070d:	ff_dbi <= 8'h04;
		14'h070e:	ff_dbi <= 8'h78;
		14'h070f:	ff_dbi <= 8'h00;
		14'h0710:	ff_dbi <= 8'h00;
		14'h0711:	ff_dbi <= 8'hfc;
		14'h0712:	ff_dbi <= 8'h02;
		14'h0713:	ff_dbi <= 8'h02;
		14'h0714:	ff_dbi <= 8'h02;
		14'h0715:	ff_dbi <= 8'h04;
		14'h0716:	ff_dbi <= 8'h18;
		14'h0717:	ff_dbi <= 8'h00;
		14'h0718:	ff_dbi <= 8'hfe;
		14'h0719:	ff_dbi <= 8'h08;
		14'h071a:	ff_dbi <= 8'h10;
		14'h071b:	ff_dbi <= 8'h20;
		14'h071c:	ff_dbi <= 8'h20;
		14'h071d:	ff_dbi <= 8'h20;
		14'h071e:	ff_dbi <= 8'h1c;
		14'h071f:	ff_dbi <= 8'h00;
		14'h0720:	ff_dbi <= 8'h20;
		14'h0721:	ff_dbi <= 8'h24;
		14'h0722:	ff_dbi <= 8'h38;
		14'h0723:	ff_dbi <= 8'h60;
		14'h0724:	ff_dbi <= 8'h80;
		14'h0725:	ff_dbi <= 8'h80;
		14'h0726:	ff_dbi <= 8'h7c;
		14'h0727:	ff_dbi <= 8'h00;
		14'h0728:	ff_dbi <= 8'h2c;
		14'h0729:	ff_dbi <= 8'hf2;
		14'h072a:	ff_dbi <= 8'h44;
		14'h072b:	ff_dbi <= 8'h44;
		14'h072c:	ff_dbi <= 8'h9c;
		14'h072d:	ff_dbi <= 8'h26;
		14'h072e:	ff_dbi <= 8'h1c;
		14'h072f:	ff_dbi <= 8'h00;
		14'h0730:	ff_dbi <= 8'h00;
		14'h0731:	ff_dbi <= 8'h9e;
		14'h0732:	ff_dbi <= 8'h80;
		14'h0733:	ff_dbi <= 8'h80;
		14'h0734:	ff_dbi <= 8'h80;
		14'h0735:	ff_dbi <= 8'h90;
		14'h0736:	ff_dbi <= 8'h4e;
		14'h0737:	ff_dbi <= 8'h00;
		14'h0738:	ff_dbi <= 8'h48;
		14'h0739:	ff_dbi <= 8'h48;
		14'h073a:	ff_dbi <= 8'h7c;
		14'h073b:	ff_dbi <= 8'hd2;
		14'h073c:	ff_dbi <= 8'hb6;
		14'h073d:	ff_dbi <= 8'haa;
		14'h073e:	ff_dbi <= 8'h4c;
		14'h073f:	ff_dbi <= 8'h00;
		14'h0740:	ff_dbi <= 8'h40;
		14'h0741:	ff_dbi <= 8'h4c;
		14'h0742:	ff_dbi <= 8'hd2;
		14'h0743:	ff_dbi <= 8'h62;
		14'h0744:	ff_dbi <= 8'h4e;
		14'h0745:	ff_dbi <= 8'hd2;
		14'h0746:	ff_dbi <= 8'h4e;
		14'h0747:	ff_dbi <= 8'h00;
		14'h0748:	ff_dbi <= 8'h00;
		14'h0749:	ff_dbi <= 8'h38;
		14'h074a:	ff_dbi <= 8'h54;
		14'h074b:	ff_dbi <= 8'h92;
		14'h074c:	ff_dbi <= 8'ha2;
		14'h074d:	ff_dbi <= 8'ha2;
		14'h074e:	ff_dbi <= 8'h44;
		14'h074f:	ff_dbi <= 8'h00;
		14'h0750:	ff_dbi <= 8'h04;
		14'h0751:	ff_dbi <= 8'h9e;
		14'h0752:	ff_dbi <= 8'h84;
		14'h0753:	ff_dbi <= 8'h84;
		14'h0754:	ff_dbi <= 8'h8c;
		14'h0755:	ff_dbi <= 8'h96;
		14'h0756:	ff_dbi <= 8'h4c;
		14'h0757:	ff_dbi <= 8'h00;
		14'h0758:	ff_dbi <= 8'h10;
		14'h0759:	ff_dbi <= 8'he4;
		14'h075a:	ff_dbi <= 8'h26;
		14'h075b:	ff_dbi <= 8'h44;
		14'h075c:	ff_dbi <= 8'h44;
		14'h075d:	ff_dbi <= 8'h48;
		14'h075e:	ff_dbi <= 8'h30;
		14'h075f:	ff_dbi <= 8'h00;
		14'h0760:	ff_dbi <= 8'h20;
		14'h0761:	ff_dbi <= 8'h10;
		14'h0762:	ff_dbi <= 8'h00;
		14'h0763:	ff_dbi <= 8'h20;
		14'h0764:	ff_dbi <= 8'h14;
		14'h0765:	ff_dbi <= 8'h52;
		14'h0766:	ff_dbi <= 8'hb2;
		14'h0767:	ff_dbi <= 8'h00;
		14'h0768:	ff_dbi <= 8'h00;
		14'h0769:	ff_dbi <= 8'h00;
		14'h076a:	ff_dbi <= 8'h20;
		14'h076b:	ff_dbi <= 8'h50;
		14'h076c:	ff_dbi <= 8'h88;
		14'h076d:	ff_dbi <= 8'h04;
		14'h076e:	ff_dbi <= 8'h02;
		14'h076f:	ff_dbi <= 8'h00;
		14'h0770:	ff_dbi <= 8'h1e;
		14'h0771:	ff_dbi <= 8'h84;
		14'h0772:	ff_dbi <= 8'h9e;
		14'h0773:	ff_dbi <= 8'h84;
		14'h0774:	ff_dbi <= 8'h8c;
		14'h0775:	ff_dbi <= 8'h96;
		14'h0776:	ff_dbi <= 8'h4c;
		14'h0777:	ff_dbi <= 8'h00;
		14'h0778:	ff_dbi <= 8'h10;
		14'h0779:	ff_dbi <= 8'hfc;
		14'h077a:	ff_dbi <= 8'h10;
		14'h077b:	ff_dbi <= 8'hfc;
		14'h077c:	ff_dbi <= 8'h70;
		14'h077d:	ff_dbi <= 8'h98;
		14'h077e:	ff_dbi <= 8'h74;
		14'h077f:	ff_dbi <= 8'h00;
		14'h0780:	ff_dbi <= 8'h70;
		14'h0781:	ff_dbi <= 8'h10;
		14'h0782:	ff_dbi <= 8'h14;
		14'h0783:	ff_dbi <= 8'h7e;
		14'h0784:	ff_dbi <= 8'ha4;
		14'h0785:	ff_dbi <= 8'ha4;
		14'h0786:	ff_dbi <= 8'h48;
		14'h0787:	ff_dbi <= 8'h00;
		14'h0788:	ff_dbi <= 8'h20;
		14'h0789:	ff_dbi <= 8'hf4;
		14'h078a:	ff_dbi <= 8'h22;
		14'h078b:	ff_dbi <= 8'h60;
		14'h078c:	ff_dbi <= 8'ha2;
		14'h078d:	ff_dbi <= 8'h62;
		14'h078e:	ff_dbi <= 8'h1c;
		14'h078f:	ff_dbi <= 8'h00;
		14'h0790:	ff_dbi <= 8'h48;
		14'h0791:	ff_dbi <= 8'h48;
		14'h0792:	ff_dbi <= 8'h7c;
		14'h0793:	ff_dbi <= 8'haa;
		14'h0794:	ff_dbi <= 8'h92;
		14'h0795:	ff_dbi <= 8'ha2;
		14'h0796:	ff_dbi <= 8'h44;
		14'h0797:	ff_dbi <= 8'h00;
		14'h0798:	ff_dbi <= 8'h20;
		14'h0799:	ff_dbi <= 8'hf8;
		14'h079a:	ff_dbi <= 8'h20;
		14'h079b:	ff_dbi <= 8'hf8;
		14'h079c:	ff_dbi <= 8'h20;
		14'h079d:	ff_dbi <= 8'h24;
		14'h079e:	ff_dbi <= 8'h18;
		14'h079f:	ff_dbi <= 8'h00;
		14'h07a0:	ff_dbi <= 8'h48;
		14'h07a1:	ff_dbi <= 8'h5c;
		14'h07a2:	ff_dbi <= 8'h6a;
		14'h07a3:	ff_dbi <= 8'he2;
		14'h07a4:	ff_dbi <= 8'h24;
		14'h07a5:	ff_dbi <= 8'h10;
		14'h07a6:	ff_dbi <= 8'h10;
		14'h07a7:	ff_dbi <= 8'h00;
		14'h07a8:	ff_dbi <= 8'h10;
		14'h07a9:	ff_dbi <= 8'h9c;
		14'h07aa:	ff_dbi <= 8'hb2;
		14'h07ab:	ff_dbi <= 8'hd2;
		14'h07ac:	ff_dbi <= 8'h92;
		14'h07ad:	ff_dbi <= 8'h1c;
		14'h07ae:	ff_dbi <= 8'h20;
		14'h07af:	ff_dbi <= 8'h00;
		14'h07b0:	ff_dbi <= 8'h10;
		14'h07b1:	ff_dbi <= 8'h1c;
		14'h07b2:	ff_dbi <= 8'h10;
		14'h07b3:	ff_dbi <= 8'h10;
		14'h07b4:	ff_dbi <= 8'h78;
		14'h07b5:	ff_dbi <= 8'h94;
		14'h07b6:	ff_dbi <= 8'h70;
		14'h07b7:	ff_dbi <= 8'h00;
		14'h07b8:	ff_dbi <= 8'h60;
		14'h07b9:	ff_dbi <= 8'h10;
		14'h07ba:	ff_dbi <= 8'h80;
		14'h07bb:	ff_dbi <= 8'hb8;
		14'h07bc:	ff_dbi <= 8'hc4;
		14'h07bd:	ff_dbi <= 8'h84;
		14'h07be:	ff_dbi <= 8'h38;
		14'h07bf:	ff_dbi <= 8'h00;
		14'h07c0:	ff_dbi <= 8'h08;
		14'h07c1:	ff_dbi <= 8'h84;
		14'h07c2:	ff_dbi <= 8'h84;
		14'h07c3:	ff_dbi <= 8'h84;
		14'h07c4:	ff_dbi <= 8'h44;
		14'h07c5:	ff_dbi <= 8'h08;
		14'h07c6:	ff_dbi <= 8'h30;
		14'h07c7:	ff_dbi <= 8'h00;
		14'h07c8:	ff_dbi <= 8'h78;
		14'h07c9:	ff_dbi <= 8'h10;
		14'h07ca:	ff_dbi <= 8'h38;
		14'h07cb:	ff_dbi <= 8'h44;
		14'h07cc:	ff_dbi <= 8'hb4;
		14'h07cd:	ff_dbi <= 8'h4c;
		14'h07ce:	ff_dbi <= 8'h38;
		14'h07cf:	ff_dbi <= 8'h00;
		14'h07d0:	ff_dbi <= 8'h20;
		14'h07d1:	ff_dbi <= 8'h2c;
		14'h07d2:	ff_dbi <= 8'hf4;
		14'h07d3:	ff_dbi <= 8'h24;
		14'h07d4:	ff_dbi <= 8'h64;
		14'h07d5:	ff_dbi <= 8'ha4;
		14'h07d6:	ff_dbi <= 8'h26;
		14'h07d7:	ff_dbi <= 8'h00;
		14'h07d8:	ff_dbi <= 8'h78;
		14'h07d9:	ff_dbi <= 8'h10;
		14'h07da:	ff_dbi <= 8'h20;
		14'h07db:	ff_dbi <= 8'h78;
		14'h07dc:	ff_dbi <= 8'h84;
		14'h07dd:	ff_dbi <= 8'h04;
		14'h07de:	ff_dbi <= 8'h38;
		14'h07df:	ff_dbi <= 8'h00;
		14'h07e0:	ff_dbi <= 8'h40;
		14'h07e1:	ff_dbi <= 8'h40;
		14'h07e2:	ff_dbi <= 8'hdc;
		14'h07e3:	ff_dbi <= 8'h62;
		14'h07e4:	ff_dbi <= 8'h42;
		14'h07e5:	ff_dbi <= 8'hc2;
		14'h07e6:	ff_dbi <= 8'h44;
		14'h07e7:	ff_dbi <= 8'h00;
		14'h07e8:	ff_dbi <= 8'h10;
		14'h07e9:	ff_dbi <= 8'h10;
		14'h07ea:	ff_dbi <= 8'h20;
		14'h07eb:	ff_dbi <= 8'h20;
		14'h07ec:	ff_dbi <= 8'h60;
		14'h07ed:	ff_dbi <= 8'h52;
		14'h07ee:	ff_dbi <= 8'h8c;
		14'h07ef:	ff_dbi <= 8'h00;
		14'h07f0:	ff_dbi <= 8'h00;
		14'h07f1:	ff_dbi <= 8'h00;
		14'h07f2:	ff_dbi <= 8'h00;
		14'h07f3:	ff_dbi <= 8'h00;
		14'h07f4:	ff_dbi <= 8'h00;
		14'h07f5:	ff_dbi <= 8'h00;
		14'h07f6:	ff_dbi <= 8'h00;
		14'h07f7:	ff_dbi <= 8'h00;
		14'h07f8:	ff_dbi <= 8'hff;
		14'h07f9:	ff_dbi <= 8'hff;
		14'h07fa:	ff_dbi <= 8'hff;
		14'h07fb:	ff_dbi <= 8'hff;
		14'h07fc:	ff_dbi <= 8'hff;
		14'h07fd:	ff_dbi <= 8'hff;
		14'h07fe:	ff_dbi <= 8'hff;
		14'h07ff:	ff_dbi <= 8'hff;
		14'h0800:	ff_dbi <= 8'h00;
		14'h0801:	ff_dbi <= 8'h00;
		14'h0802:	ff_dbi <= 8'h00;
		14'h0803:	ff_dbi <= 8'h00;
		14'h0804:	ff_dbi <= 8'h00;
		14'h0805:	ff_dbi <= 8'h00;
		14'h0806:	ff_dbi <= 8'h00;
		14'h0807:	ff_dbi <= 8'h00;
		14'h0808:	ff_dbi <= 8'h00;
		14'h0809:	ff_dbi <= 8'h00;
		14'h080a:	ff_dbi <= 8'h00;
		14'h080b:	ff_dbi <= 8'h00;
		14'h080c:	ff_dbi <= 8'h00;
		14'h080d:	ff_dbi <= 8'h00;
		14'h080e:	ff_dbi <= 8'h00;
		14'h080f:	ff_dbi <= 8'h00;
		14'h0810:	ff_dbi <= 8'h00;
		14'h0811:	ff_dbi <= 8'h00;
		14'h0812:	ff_dbi <= 8'h00;
		14'h0813:	ff_dbi <= 8'h00;
		14'h0814:	ff_dbi <= 8'h00;
		14'h0815:	ff_dbi <= 8'h00;
		14'h0816:	ff_dbi <= 8'h00;
		14'h0817:	ff_dbi <= 8'h00;
		14'h0818:	ff_dbi <= 8'h00;
		14'h0819:	ff_dbi <= 8'h00;
		14'h081a:	ff_dbi <= 8'h00;
		14'h081b:	ff_dbi <= 8'h00;
		14'h081c:	ff_dbi <= 8'h00;
		14'h081d:	ff_dbi <= 8'h00;
		14'h081e:	ff_dbi <= 8'h00;
		14'h081f:	ff_dbi <= 8'h00;
		14'h0820:	ff_dbi <= 8'h00;
		14'h0821:	ff_dbi <= 8'h00;
		14'h0822:	ff_dbi <= 8'h00;
		14'h0823:	ff_dbi <= 8'h00;
		14'h0824:	ff_dbi <= 8'h00;
		14'h0825:	ff_dbi <= 8'h00;
		14'h0826:	ff_dbi <= 8'h00;
		14'h0827:	ff_dbi <= 8'h00;
		14'h0828:	ff_dbi <= 8'h00;
		14'h0829:	ff_dbi <= 8'h00;
		14'h082a:	ff_dbi <= 8'h00;
		14'h082b:	ff_dbi <= 8'h00;
		14'h082c:	ff_dbi <= 8'h00;
		14'h082d:	ff_dbi <= 8'h00;
		14'h082e:	ff_dbi <= 8'h00;
		14'h082f:	ff_dbi <= 8'h00;
		14'h0830:	ff_dbi <= 8'h00;
		14'h0831:	ff_dbi <= 8'h00;
		14'h0832:	ff_dbi <= 8'h00;
		14'h0833:	ff_dbi <= 8'h00;
		14'h0834:	ff_dbi <= 8'h00;
		14'h0835:	ff_dbi <= 8'h00;
		14'h0836:	ff_dbi <= 8'h00;
		14'h0837:	ff_dbi <= 8'h00;
		14'h0838:	ff_dbi <= 8'h00;
		14'h0839:	ff_dbi <= 8'h00;
		14'h083a:	ff_dbi <= 8'h00;
		14'h083b:	ff_dbi <= 8'h00;
		14'h083c:	ff_dbi <= 8'h00;
		14'h083d:	ff_dbi <= 8'h00;
		14'h083e:	ff_dbi <= 8'h00;
		14'h083f:	ff_dbi <= 8'h00;
		14'h0840:	ff_dbi <= 8'h00;
		14'h0841:	ff_dbi <= 8'h00;
		14'h0842:	ff_dbi <= 8'h00;
		14'h0843:	ff_dbi <= 8'h00;
		14'h0844:	ff_dbi <= 8'h00;
		14'h0845:	ff_dbi <= 8'h00;
		14'h0846:	ff_dbi <= 8'h00;
		14'h0847:	ff_dbi <= 8'h00;
		14'h0848:	ff_dbi <= 8'h00;
		14'h0849:	ff_dbi <= 8'h00;
		14'h084a:	ff_dbi <= 8'h00;
		14'h084b:	ff_dbi <= 8'h00;
		14'h084c:	ff_dbi <= 8'h00;
		14'h084d:	ff_dbi <= 8'h00;
		14'h084e:	ff_dbi <= 8'h00;
		14'h084f:	ff_dbi <= 8'h00;
		14'h0850:	ff_dbi <= 8'h00;
		14'h0851:	ff_dbi <= 8'h00;
		14'h0852:	ff_dbi <= 8'h00;
		14'h0853:	ff_dbi <= 8'h00;
		14'h0854:	ff_dbi <= 8'h00;
		14'h0855:	ff_dbi <= 8'h00;
		14'h0856:	ff_dbi <= 8'h00;
		14'h0857:	ff_dbi <= 8'h00;
		14'h0858:	ff_dbi <= 8'h00;
		14'h0859:	ff_dbi <= 8'h00;
		14'h085a:	ff_dbi <= 8'h00;
		14'h085b:	ff_dbi <= 8'h00;
		14'h085c:	ff_dbi <= 8'h00;
		14'h085d:	ff_dbi <= 8'h00;
		14'h085e:	ff_dbi <= 8'h00;
		14'h085f:	ff_dbi <= 8'h00;
		14'h0860:	ff_dbi <= 8'h00;
		14'h0861:	ff_dbi <= 8'h00;
		14'h0862:	ff_dbi <= 8'h00;
		14'h0863:	ff_dbi <= 8'h00;
		14'h0864:	ff_dbi <= 8'h00;
		14'h0865:	ff_dbi <= 8'h00;
		14'h0866:	ff_dbi <= 8'h00;
		14'h0867:	ff_dbi <= 8'h00;
		14'h0868:	ff_dbi <= 8'h00;
		14'h0869:	ff_dbi <= 8'h00;
		14'h086a:	ff_dbi <= 8'h00;
		14'h086b:	ff_dbi <= 8'h00;
		14'h086c:	ff_dbi <= 8'h00;
		14'h086d:	ff_dbi <= 8'h00;
		14'h086e:	ff_dbi <= 8'h00;
		14'h086f:	ff_dbi <= 8'h00;
		14'h0870:	ff_dbi <= 8'h00;
		14'h0871:	ff_dbi <= 8'h00;
		14'h0872:	ff_dbi <= 8'h00;
		14'h0873:	ff_dbi <= 8'h00;
		14'h0874:	ff_dbi <= 8'h00;
		14'h0875:	ff_dbi <= 8'h00;
		14'h0876:	ff_dbi <= 8'h00;
		14'h0877:	ff_dbi <= 8'h00;
		14'h0878:	ff_dbi <= 8'h00;
		14'h0879:	ff_dbi <= 8'h00;
		14'h087a:	ff_dbi <= 8'h00;
		14'h087b:	ff_dbi <= 8'h00;
		14'h087c:	ff_dbi <= 8'h00;
		14'h087d:	ff_dbi <= 8'h00;
		14'h087e:	ff_dbi <= 8'h00;
		14'h087f:	ff_dbi <= 8'h00;
		14'h0880:	ff_dbi <= 8'h00;
		14'h0881:	ff_dbi <= 8'h00;
		14'h0882:	ff_dbi <= 8'h00;
		14'h0883:	ff_dbi <= 8'h00;
		14'h0884:	ff_dbi <= 8'h00;
		14'h0885:	ff_dbi <= 8'h00;
		14'h0886:	ff_dbi <= 8'h00;
		14'h0887:	ff_dbi <= 8'h00;
		14'h0888:	ff_dbi <= 8'h00;
		14'h0889:	ff_dbi <= 8'h00;
		14'h088a:	ff_dbi <= 8'h00;
		14'h088b:	ff_dbi <= 8'h00;
		14'h088c:	ff_dbi <= 8'h00;
		14'h088d:	ff_dbi <= 8'h00;
		14'h088e:	ff_dbi <= 8'h00;
		14'h088f:	ff_dbi <= 8'h00;
		14'h0890:	ff_dbi <= 8'h00;
		14'h0891:	ff_dbi <= 8'h00;
		14'h0892:	ff_dbi <= 8'h00;
		14'h0893:	ff_dbi <= 8'h00;
		14'h0894:	ff_dbi <= 8'h00;
		14'h0895:	ff_dbi <= 8'h00;
		14'h0896:	ff_dbi <= 8'h00;
		14'h0897:	ff_dbi <= 8'h00;
		14'h0898:	ff_dbi <= 8'h00;
		14'h0899:	ff_dbi <= 8'h00;
		14'h089a:	ff_dbi <= 8'h00;
		14'h089b:	ff_dbi <= 8'h00;
		14'h089c:	ff_dbi <= 8'h00;
		14'h089d:	ff_dbi <= 8'h00;
		14'h089e:	ff_dbi <= 8'h00;
		14'h089f:	ff_dbi <= 8'h00;
		14'h08a0:	ff_dbi <= 8'h00;
		14'h08a1:	ff_dbi <= 8'h00;
		14'h08a2:	ff_dbi <= 8'h00;
		14'h08a3:	ff_dbi <= 8'h00;
		14'h08a4:	ff_dbi <= 8'h00;
		14'h08a5:	ff_dbi <= 8'h00;
		14'h08a6:	ff_dbi <= 8'h00;
		14'h08a7:	ff_dbi <= 8'h00;
		14'h08a8:	ff_dbi <= 8'h00;
		14'h08a9:	ff_dbi <= 8'h00;
		14'h08aa:	ff_dbi <= 8'h00;
		14'h08ab:	ff_dbi <= 8'h00;
		14'h08ac:	ff_dbi <= 8'h00;
		14'h08ad:	ff_dbi <= 8'h00;
		14'h08ae:	ff_dbi <= 8'h00;
		14'h08af:	ff_dbi <= 8'h00;
		14'h08b0:	ff_dbi <= 8'h00;
		14'h08b1:	ff_dbi <= 8'h00;
		14'h08b2:	ff_dbi <= 8'h00;
		14'h08b3:	ff_dbi <= 8'h00;
		14'h08b4:	ff_dbi <= 8'h00;
		14'h08b5:	ff_dbi <= 8'h00;
		14'h08b6:	ff_dbi <= 8'h00;
		14'h08b7:	ff_dbi <= 8'h00;
		14'h08b8:	ff_dbi <= 8'h00;
		14'h08b9:	ff_dbi <= 8'h00;
		14'h08ba:	ff_dbi <= 8'h00;
		14'h08bb:	ff_dbi <= 8'h00;
		14'h08bc:	ff_dbi <= 8'h00;
		14'h08bd:	ff_dbi <= 8'h00;
		14'h08be:	ff_dbi <= 8'h00;
		14'h08bf:	ff_dbi <= 8'h00;
		14'h08c0:	ff_dbi <= 8'h00;
		14'h08c1:	ff_dbi <= 8'h00;
		14'h08c2:	ff_dbi <= 8'h00;
		14'h08c3:	ff_dbi <= 8'h00;
		14'h08c4:	ff_dbi <= 8'h00;
		14'h08c5:	ff_dbi <= 8'h00;
		14'h08c6:	ff_dbi <= 8'h00;
		14'h08c7:	ff_dbi <= 8'h00;
		14'h08c8:	ff_dbi <= 8'h00;
		14'h08c9:	ff_dbi <= 8'h00;
		14'h08ca:	ff_dbi <= 8'h00;
		14'h08cb:	ff_dbi <= 8'h00;
		14'h08cc:	ff_dbi <= 8'h00;
		14'h08cd:	ff_dbi <= 8'h00;
		14'h08ce:	ff_dbi <= 8'h00;
		14'h08cf:	ff_dbi <= 8'h00;
		14'h08d0:	ff_dbi <= 8'h00;
		14'h08d1:	ff_dbi <= 8'h00;
		14'h08d2:	ff_dbi <= 8'h00;
		14'h08d3:	ff_dbi <= 8'h00;
		14'h08d4:	ff_dbi <= 8'h00;
		14'h08d5:	ff_dbi <= 8'h00;
		14'h08d6:	ff_dbi <= 8'h00;
		14'h08d7:	ff_dbi <= 8'h00;
		14'h08d8:	ff_dbi <= 8'h00;
		14'h08d9:	ff_dbi <= 8'h00;
		14'h08da:	ff_dbi <= 8'h00;
		14'h08db:	ff_dbi <= 8'h00;
		14'h08dc:	ff_dbi <= 8'h00;
		14'h08dd:	ff_dbi <= 8'h00;
		14'h08de:	ff_dbi <= 8'h00;
		14'h08df:	ff_dbi <= 8'h00;
		14'h08e0:	ff_dbi <= 8'h00;
		14'h08e1:	ff_dbi <= 8'h00;
		14'h08e2:	ff_dbi <= 8'h00;
		14'h08e3:	ff_dbi <= 8'h00;
		14'h08e4:	ff_dbi <= 8'h00;
		14'h08e5:	ff_dbi <= 8'h00;
		14'h08e6:	ff_dbi <= 8'h00;
		14'h08e7:	ff_dbi <= 8'h00;
		14'h08e8:	ff_dbi <= 8'h00;
		14'h08e9:	ff_dbi <= 8'h00;
		14'h08ea:	ff_dbi <= 8'h00;
		14'h08eb:	ff_dbi <= 8'h00;
		14'h08ec:	ff_dbi <= 8'h00;
		14'h08ed:	ff_dbi <= 8'h00;
		14'h08ee:	ff_dbi <= 8'h00;
		14'h08ef:	ff_dbi <= 8'h00;
		14'h08f0:	ff_dbi <= 8'h00;
		14'h08f1:	ff_dbi <= 8'h00;
		14'h08f2:	ff_dbi <= 8'h00;
		14'h08f3:	ff_dbi <= 8'h00;
		14'h08f4:	ff_dbi <= 8'h00;
		14'h08f5:	ff_dbi <= 8'h00;
		14'h08f6:	ff_dbi <= 8'h00;
		14'h08f7:	ff_dbi <= 8'h00;
		14'h08f8:	ff_dbi <= 8'h00;
		14'h08f9:	ff_dbi <= 8'h00;
		14'h08fa:	ff_dbi <= 8'h00;
		14'h08fb:	ff_dbi <= 8'h00;
		14'h08fc:	ff_dbi <= 8'h00;
		14'h08fd:	ff_dbi <= 8'h00;
		14'h08fe:	ff_dbi <= 8'h00;
		14'h08ff:	ff_dbi <= 8'h00;
		14'h0900:	ff_dbi <= 8'h00;
		14'h0901:	ff_dbi <= 8'h00;
		14'h0902:	ff_dbi <= 8'h00;
		14'h0903:	ff_dbi <= 8'h00;
		14'h0904:	ff_dbi <= 8'h00;
		14'h0905:	ff_dbi <= 8'h00;
		14'h0906:	ff_dbi <= 8'h00;
		14'h0907:	ff_dbi <= 8'h00;
		14'h0908:	ff_dbi <= 8'h00;
		14'h0909:	ff_dbi <= 8'h00;
		14'h090a:	ff_dbi <= 8'h00;
		14'h090b:	ff_dbi <= 8'h00;
		14'h090c:	ff_dbi <= 8'h00;
		14'h090d:	ff_dbi <= 8'h00;
		14'h090e:	ff_dbi <= 8'h00;
		14'h090f:	ff_dbi <= 8'h00;
		14'h0910:	ff_dbi <= 8'h00;
		14'h0911:	ff_dbi <= 8'h00;
		14'h0912:	ff_dbi <= 8'h00;
		14'h0913:	ff_dbi <= 8'h00;
		14'h0914:	ff_dbi <= 8'h00;
		14'h0915:	ff_dbi <= 8'h00;
		14'h0916:	ff_dbi <= 8'h00;
		14'h0917:	ff_dbi <= 8'h00;
		14'h0918:	ff_dbi <= 8'h00;
		14'h0919:	ff_dbi <= 8'h00;
		14'h091a:	ff_dbi <= 8'h00;
		14'h091b:	ff_dbi <= 8'h00;
		14'h091c:	ff_dbi <= 8'h00;
		14'h091d:	ff_dbi <= 8'h00;
		14'h091e:	ff_dbi <= 8'h00;
		14'h091f:	ff_dbi <= 8'h00;
		14'h0920:	ff_dbi <= 8'h00;
		14'h0921:	ff_dbi <= 8'h00;
		14'h0922:	ff_dbi <= 8'h00;
		14'h0923:	ff_dbi <= 8'h00;
		14'h0924:	ff_dbi <= 8'h00;
		14'h0925:	ff_dbi <= 8'h00;
		14'h0926:	ff_dbi <= 8'h00;
		14'h0927:	ff_dbi <= 8'h00;
		14'h0928:	ff_dbi <= 8'h00;
		14'h0929:	ff_dbi <= 8'h00;
		14'h092a:	ff_dbi <= 8'h00;
		14'h092b:	ff_dbi <= 8'h00;
		14'h092c:	ff_dbi <= 8'h00;
		14'h092d:	ff_dbi <= 8'h00;
		14'h092e:	ff_dbi <= 8'h00;
		14'h092f:	ff_dbi <= 8'h00;
		14'h0930:	ff_dbi <= 8'h00;
		14'h0931:	ff_dbi <= 8'h00;
		14'h0932:	ff_dbi <= 8'h00;
		14'h0933:	ff_dbi <= 8'h00;
		14'h0934:	ff_dbi <= 8'h00;
		14'h0935:	ff_dbi <= 8'h00;
		14'h0936:	ff_dbi <= 8'h00;
		14'h0937:	ff_dbi <= 8'h00;
		14'h0938:	ff_dbi <= 8'h00;
		14'h0939:	ff_dbi <= 8'h00;
		14'h093a:	ff_dbi <= 8'h00;
		14'h093b:	ff_dbi <= 8'h00;
		14'h093c:	ff_dbi <= 8'h00;
		14'h093d:	ff_dbi <= 8'h00;
		14'h093e:	ff_dbi <= 8'h00;
		14'h093f:	ff_dbi <= 8'h00;
		14'h0940:	ff_dbi <= 8'h00;
		14'h0941:	ff_dbi <= 8'h00;
		14'h0942:	ff_dbi <= 8'h00;
		14'h0943:	ff_dbi <= 8'h00;
		14'h0944:	ff_dbi <= 8'h00;
		14'h0945:	ff_dbi <= 8'h00;
		14'h0946:	ff_dbi <= 8'h00;
		14'h0947:	ff_dbi <= 8'h00;
		14'h0948:	ff_dbi <= 8'h00;
		14'h0949:	ff_dbi <= 8'h00;
		14'h094a:	ff_dbi <= 8'h00;
		14'h094b:	ff_dbi <= 8'h00;
		14'h094c:	ff_dbi <= 8'h00;
		14'h094d:	ff_dbi <= 8'h00;
		14'h094e:	ff_dbi <= 8'h00;
		14'h094f:	ff_dbi <= 8'h00;
		14'h0950:	ff_dbi <= 8'h00;
		14'h0951:	ff_dbi <= 8'h00;
		14'h0952:	ff_dbi <= 8'h00;
		14'h0953:	ff_dbi <= 8'h00;
		14'h0954:	ff_dbi <= 8'h00;
		14'h0955:	ff_dbi <= 8'h00;
		14'h0956:	ff_dbi <= 8'h00;
		14'h0957:	ff_dbi <= 8'h00;
		14'h0958:	ff_dbi <= 8'h00;
		14'h0959:	ff_dbi <= 8'h00;
		14'h095a:	ff_dbi <= 8'h00;
		14'h095b:	ff_dbi <= 8'h00;
		14'h095c:	ff_dbi <= 8'h00;
		14'h095d:	ff_dbi <= 8'h00;
		14'h095e:	ff_dbi <= 8'h00;
		14'h095f:	ff_dbi <= 8'h00;
		14'h0960:	ff_dbi <= 8'h00;
		14'h0961:	ff_dbi <= 8'h00;
		14'h0962:	ff_dbi <= 8'h00;
		14'h0963:	ff_dbi <= 8'h00;
		14'h0964:	ff_dbi <= 8'h00;
		14'h0965:	ff_dbi <= 8'h00;
		14'h0966:	ff_dbi <= 8'h00;
		14'h0967:	ff_dbi <= 8'h00;
		14'h0968:	ff_dbi <= 8'h00;
		14'h0969:	ff_dbi <= 8'h00;
		14'h096a:	ff_dbi <= 8'h00;
		14'h096b:	ff_dbi <= 8'h00;
		14'h096c:	ff_dbi <= 8'h00;
		14'h096d:	ff_dbi <= 8'h00;
		14'h096e:	ff_dbi <= 8'h00;
		14'h096f:	ff_dbi <= 8'h00;
		14'h0970:	ff_dbi <= 8'h00;
		14'h0971:	ff_dbi <= 8'h00;
		14'h0972:	ff_dbi <= 8'h00;
		14'h0973:	ff_dbi <= 8'h00;
		14'h0974:	ff_dbi <= 8'h00;
		14'h0975:	ff_dbi <= 8'h00;
		14'h0976:	ff_dbi <= 8'h00;
		14'h0977:	ff_dbi <= 8'h00;
		14'h0978:	ff_dbi <= 8'h00;
		14'h0979:	ff_dbi <= 8'h00;
		14'h097a:	ff_dbi <= 8'h00;
		14'h097b:	ff_dbi <= 8'h00;
		14'h097c:	ff_dbi <= 8'h00;
		14'h097d:	ff_dbi <= 8'h00;
		14'h097e:	ff_dbi <= 8'h00;
		14'h097f:	ff_dbi <= 8'h00;
		14'h0980:	ff_dbi <= 8'h00;
		14'h0981:	ff_dbi <= 8'h00;
		14'h0982:	ff_dbi <= 8'h00;
		14'h0983:	ff_dbi <= 8'h00;
		14'h0984:	ff_dbi <= 8'h00;
		14'h0985:	ff_dbi <= 8'h00;
		14'h0986:	ff_dbi <= 8'h00;
		14'h0987:	ff_dbi <= 8'h00;
		14'h0988:	ff_dbi <= 8'h00;
		14'h0989:	ff_dbi <= 8'h00;
		14'h098a:	ff_dbi <= 8'h00;
		14'h098b:	ff_dbi <= 8'h00;
		14'h098c:	ff_dbi <= 8'h00;
		14'h098d:	ff_dbi <= 8'h00;
		14'h098e:	ff_dbi <= 8'h00;
		14'h098f:	ff_dbi <= 8'h00;
		14'h0990:	ff_dbi <= 8'h00;
		14'h0991:	ff_dbi <= 8'h00;
		14'h0992:	ff_dbi <= 8'h00;
		14'h0993:	ff_dbi <= 8'h00;
		14'h0994:	ff_dbi <= 8'h00;
		14'h0995:	ff_dbi <= 8'h00;
		14'h0996:	ff_dbi <= 8'h00;
		14'h0997:	ff_dbi <= 8'h00;
		14'h0998:	ff_dbi <= 8'h00;
		14'h0999:	ff_dbi <= 8'h00;
		14'h099a:	ff_dbi <= 8'h00;
		14'h099b:	ff_dbi <= 8'h00;
		14'h099c:	ff_dbi <= 8'h00;
		14'h099d:	ff_dbi <= 8'h00;
		14'h099e:	ff_dbi <= 8'h00;
		14'h099f:	ff_dbi <= 8'h00;
		14'h09a0:	ff_dbi <= 8'h00;
		14'h09a1:	ff_dbi <= 8'h00;
		14'h09a2:	ff_dbi <= 8'h00;
		14'h09a3:	ff_dbi <= 8'h00;
		14'h09a4:	ff_dbi <= 8'h00;
		14'h09a5:	ff_dbi <= 8'h00;
		14'h09a6:	ff_dbi <= 8'h00;
		14'h09a7:	ff_dbi <= 8'h00;
		14'h09a8:	ff_dbi <= 8'h00;
		14'h09a9:	ff_dbi <= 8'h00;
		14'h09aa:	ff_dbi <= 8'h00;
		14'h09ab:	ff_dbi <= 8'h00;
		14'h09ac:	ff_dbi <= 8'h00;
		14'h09ad:	ff_dbi <= 8'h00;
		14'h09ae:	ff_dbi <= 8'h00;
		14'h09af:	ff_dbi <= 8'h00;
		14'h09b0:	ff_dbi <= 8'h00;
		14'h09b1:	ff_dbi <= 8'h00;
		14'h09b2:	ff_dbi <= 8'h00;
		14'h09b3:	ff_dbi <= 8'h00;
		14'h09b4:	ff_dbi <= 8'h00;
		14'h09b5:	ff_dbi <= 8'h00;
		14'h09b6:	ff_dbi <= 8'h00;
		14'h09b7:	ff_dbi <= 8'h00;
		14'h09b8:	ff_dbi <= 8'h00;
		14'h09b9:	ff_dbi <= 8'h00;
		14'h09ba:	ff_dbi <= 8'h00;
		14'h09bb:	ff_dbi <= 8'h00;
		14'h09bc:	ff_dbi <= 8'h00;
		14'h09bd:	ff_dbi <= 8'h00;
		14'h09be:	ff_dbi <= 8'h00;
		14'h09bf:	ff_dbi <= 8'h00;
		14'h09c0:	ff_dbi <= 8'h00;
		14'h09c1:	ff_dbi <= 8'h00;
		14'h09c2:	ff_dbi <= 8'h00;
		14'h09c3:	ff_dbi <= 8'h00;
		14'h09c4:	ff_dbi <= 8'h00;
		14'h09c5:	ff_dbi <= 8'h00;
		14'h09c6:	ff_dbi <= 8'h00;
		14'h09c7:	ff_dbi <= 8'h00;
		14'h09c8:	ff_dbi <= 8'h00;
		14'h09c9:	ff_dbi <= 8'h00;
		14'h09ca:	ff_dbi <= 8'h00;
		14'h09cb:	ff_dbi <= 8'h00;
		14'h09cc:	ff_dbi <= 8'h00;
		14'h09cd:	ff_dbi <= 8'h00;
		14'h09ce:	ff_dbi <= 8'h00;
		14'h09cf:	ff_dbi <= 8'h00;
		14'h09d0:	ff_dbi <= 8'h00;
		14'h09d1:	ff_dbi <= 8'h00;
		14'h09d2:	ff_dbi <= 8'h00;
		14'h09d3:	ff_dbi <= 8'h00;
		14'h09d4:	ff_dbi <= 8'h00;
		14'h09d5:	ff_dbi <= 8'h00;
		14'h09d6:	ff_dbi <= 8'h00;
		14'h09d7:	ff_dbi <= 8'h00;
		14'h09d8:	ff_dbi <= 8'h00;
		14'h09d9:	ff_dbi <= 8'h00;
		14'h09da:	ff_dbi <= 8'h00;
		14'h09db:	ff_dbi <= 8'h00;
		14'h09dc:	ff_dbi <= 8'h00;
		14'h09dd:	ff_dbi <= 8'h00;
		14'h09de:	ff_dbi <= 8'h00;
		14'h09df:	ff_dbi <= 8'h00;
		14'h09e0:	ff_dbi <= 8'h00;
		14'h09e1:	ff_dbi <= 8'h00;
		14'h09e2:	ff_dbi <= 8'h00;
		14'h09e3:	ff_dbi <= 8'h00;
		14'h09e4:	ff_dbi <= 8'h00;
		14'h09e5:	ff_dbi <= 8'h00;
		14'h09e6:	ff_dbi <= 8'h00;
		14'h09e7:	ff_dbi <= 8'h00;
		14'h09e8:	ff_dbi <= 8'h00;
		14'h09e9:	ff_dbi <= 8'h00;
		14'h09ea:	ff_dbi <= 8'h00;
		14'h09eb:	ff_dbi <= 8'h00;
		14'h09ec:	ff_dbi <= 8'h00;
		14'h09ed:	ff_dbi <= 8'h00;
		14'h09ee:	ff_dbi <= 8'h00;
		14'h09ef:	ff_dbi <= 8'h00;
		14'h09f0:	ff_dbi <= 8'h00;
		14'h09f1:	ff_dbi <= 8'h00;
		14'h09f2:	ff_dbi <= 8'h00;
		14'h09f3:	ff_dbi <= 8'h00;
		14'h09f4:	ff_dbi <= 8'h00;
		14'h09f5:	ff_dbi <= 8'h00;
		14'h09f6:	ff_dbi <= 8'h00;
		14'h09f7:	ff_dbi <= 8'h00;
		14'h09f8:	ff_dbi <= 8'h00;
		14'h09f9:	ff_dbi <= 8'h00;
		14'h09fa:	ff_dbi <= 8'h00;
		14'h09fb:	ff_dbi <= 8'h00;
		14'h09fc:	ff_dbi <= 8'h00;
		14'h09fd:	ff_dbi <= 8'h00;
		14'h09fe:	ff_dbi <= 8'h00;
		14'h09ff:	ff_dbi <= 8'h00;
		14'h0a00:	ff_dbi <= 8'h00;
		14'h0a01:	ff_dbi <= 8'h00;
		14'h0a02:	ff_dbi <= 8'h00;
		14'h0a03:	ff_dbi <= 8'h00;
		14'h0a04:	ff_dbi <= 8'h00;
		14'h0a05:	ff_dbi <= 8'h00;
		14'h0a06:	ff_dbi <= 8'h00;
		14'h0a07:	ff_dbi <= 8'h00;
		14'h0a08:	ff_dbi <= 8'h00;
		14'h0a09:	ff_dbi <= 8'h00;
		14'h0a0a:	ff_dbi <= 8'h00;
		14'h0a0b:	ff_dbi <= 8'h00;
		14'h0a0c:	ff_dbi <= 8'h00;
		14'h0a0d:	ff_dbi <= 8'h00;
		14'h0a0e:	ff_dbi <= 8'h00;
		14'h0a0f:	ff_dbi <= 8'h00;
		14'h0a10:	ff_dbi <= 8'h00;
		14'h0a11:	ff_dbi <= 8'h00;
		14'h0a12:	ff_dbi <= 8'h00;
		14'h0a13:	ff_dbi <= 8'h00;
		14'h0a14:	ff_dbi <= 8'h00;
		14'h0a15:	ff_dbi <= 8'h00;
		14'h0a16:	ff_dbi <= 8'h00;
		14'h0a17:	ff_dbi <= 8'h00;
		14'h0a18:	ff_dbi <= 8'h00;
		14'h0a19:	ff_dbi <= 8'h00;
		14'h0a1a:	ff_dbi <= 8'h00;
		14'h0a1b:	ff_dbi <= 8'h00;
		14'h0a1c:	ff_dbi <= 8'h00;
		14'h0a1d:	ff_dbi <= 8'h00;
		14'h0a1e:	ff_dbi <= 8'h00;
		14'h0a1f:	ff_dbi <= 8'h00;
		14'h0a20:	ff_dbi <= 8'h00;
		14'h0a21:	ff_dbi <= 8'h00;
		14'h0a22:	ff_dbi <= 8'h00;
		14'h0a23:	ff_dbi <= 8'h00;
		14'h0a24:	ff_dbi <= 8'h00;
		14'h0a25:	ff_dbi <= 8'h00;
		14'h0a26:	ff_dbi <= 8'h00;
		14'h0a27:	ff_dbi <= 8'h00;
		14'h0a28:	ff_dbi <= 8'h00;
		14'h0a29:	ff_dbi <= 8'h00;
		14'h0a2a:	ff_dbi <= 8'h00;
		14'h0a2b:	ff_dbi <= 8'h00;
		14'h0a2c:	ff_dbi <= 8'h00;
		14'h0a2d:	ff_dbi <= 8'h00;
		14'h0a2e:	ff_dbi <= 8'h00;
		14'h0a2f:	ff_dbi <= 8'h00;
		14'h0a30:	ff_dbi <= 8'h00;
		14'h0a31:	ff_dbi <= 8'h00;
		14'h0a32:	ff_dbi <= 8'h00;
		14'h0a33:	ff_dbi <= 8'h00;
		14'h0a34:	ff_dbi <= 8'h00;
		14'h0a35:	ff_dbi <= 8'h00;
		14'h0a36:	ff_dbi <= 8'h00;
		14'h0a37:	ff_dbi <= 8'h00;
		14'h0a38:	ff_dbi <= 8'h00;
		14'h0a39:	ff_dbi <= 8'h00;
		14'h0a3a:	ff_dbi <= 8'h00;
		14'h0a3b:	ff_dbi <= 8'h00;
		14'h0a3c:	ff_dbi <= 8'h00;
		14'h0a3d:	ff_dbi <= 8'h00;
		14'h0a3e:	ff_dbi <= 8'h00;
		14'h0a3f:	ff_dbi <= 8'h00;
		14'h0a40:	ff_dbi <= 8'h00;
		14'h0a41:	ff_dbi <= 8'h00;
		14'h0a42:	ff_dbi <= 8'h00;
		14'h0a43:	ff_dbi <= 8'h00;
		14'h0a44:	ff_dbi <= 8'h00;
		14'h0a45:	ff_dbi <= 8'h00;
		14'h0a46:	ff_dbi <= 8'h00;
		14'h0a47:	ff_dbi <= 8'h00;
		14'h0a48:	ff_dbi <= 8'h00;
		14'h0a49:	ff_dbi <= 8'h00;
		14'h0a4a:	ff_dbi <= 8'h00;
		14'h0a4b:	ff_dbi <= 8'h00;
		14'h0a4c:	ff_dbi <= 8'h00;
		14'h0a4d:	ff_dbi <= 8'h00;
		14'h0a4e:	ff_dbi <= 8'h00;
		14'h0a4f:	ff_dbi <= 8'h00;
		14'h0a50:	ff_dbi <= 8'h00;
		14'h0a51:	ff_dbi <= 8'h00;
		14'h0a52:	ff_dbi <= 8'h00;
		14'h0a53:	ff_dbi <= 8'h00;
		14'h0a54:	ff_dbi <= 8'h00;
		14'h0a55:	ff_dbi <= 8'h00;
		14'h0a56:	ff_dbi <= 8'h00;
		14'h0a57:	ff_dbi <= 8'h00;
		14'h0a58:	ff_dbi <= 8'h00;
		14'h0a59:	ff_dbi <= 8'h00;
		14'h0a5a:	ff_dbi <= 8'h00;
		14'h0a5b:	ff_dbi <= 8'h00;
		14'h0a5c:	ff_dbi <= 8'h00;
		14'h0a5d:	ff_dbi <= 8'h00;
		14'h0a5e:	ff_dbi <= 8'h00;
		14'h0a5f:	ff_dbi <= 8'h00;
		14'h0a60:	ff_dbi <= 8'h00;
		14'h0a61:	ff_dbi <= 8'h00;
		14'h0a62:	ff_dbi <= 8'h00;
		14'h0a63:	ff_dbi <= 8'h00;
		14'h0a64:	ff_dbi <= 8'h00;
		14'h0a65:	ff_dbi <= 8'h00;
		14'h0a66:	ff_dbi <= 8'h00;
		14'h0a67:	ff_dbi <= 8'h00;
		14'h0a68:	ff_dbi <= 8'h00;
		14'h0a69:	ff_dbi <= 8'h00;
		14'h0a6a:	ff_dbi <= 8'h00;
		14'h0a6b:	ff_dbi <= 8'h00;
		14'h0a6c:	ff_dbi <= 8'h00;
		14'h0a6d:	ff_dbi <= 8'h00;
		14'h0a6e:	ff_dbi <= 8'h00;
		14'h0a6f:	ff_dbi <= 8'h00;
		14'h0a70:	ff_dbi <= 8'h00;
		14'h0a71:	ff_dbi <= 8'h00;
		14'h0a72:	ff_dbi <= 8'h00;
		14'h0a73:	ff_dbi <= 8'h00;
		14'h0a74:	ff_dbi <= 8'h00;
		14'h0a75:	ff_dbi <= 8'h00;
		14'h0a76:	ff_dbi <= 8'h00;
		14'h0a77:	ff_dbi <= 8'h00;
		14'h0a78:	ff_dbi <= 8'h00;
		14'h0a79:	ff_dbi <= 8'h00;
		14'h0a7a:	ff_dbi <= 8'h00;
		14'h0a7b:	ff_dbi <= 8'h00;
		14'h0a7c:	ff_dbi <= 8'h00;
		14'h0a7d:	ff_dbi <= 8'h00;
		14'h0a7e:	ff_dbi <= 8'h00;
		14'h0a7f:	ff_dbi <= 8'h00;
		14'h0a80:	ff_dbi <= 8'h00;
		14'h0a81:	ff_dbi <= 8'h00;
		14'h0a82:	ff_dbi <= 8'h00;
		14'h0a83:	ff_dbi <= 8'h00;
		14'h0a84:	ff_dbi <= 8'h00;
		14'h0a85:	ff_dbi <= 8'h00;
		14'h0a86:	ff_dbi <= 8'h00;
		14'h0a87:	ff_dbi <= 8'h00;
		14'h0a88:	ff_dbi <= 8'h00;
		14'h0a89:	ff_dbi <= 8'h00;
		14'h0a8a:	ff_dbi <= 8'h00;
		14'h0a8b:	ff_dbi <= 8'h00;
		14'h0a8c:	ff_dbi <= 8'h00;
		14'h0a8d:	ff_dbi <= 8'h00;
		14'h0a8e:	ff_dbi <= 8'h00;
		14'h0a8f:	ff_dbi <= 8'h00;
		14'h0a90:	ff_dbi <= 8'h00;
		14'h0a91:	ff_dbi <= 8'h00;
		14'h0a92:	ff_dbi <= 8'h00;
		14'h0a93:	ff_dbi <= 8'h00;
		14'h0a94:	ff_dbi <= 8'h00;
		14'h0a95:	ff_dbi <= 8'h00;
		14'h0a96:	ff_dbi <= 8'h00;
		14'h0a97:	ff_dbi <= 8'h00;
		14'h0a98:	ff_dbi <= 8'h00;
		14'h0a99:	ff_dbi <= 8'h00;
		14'h0a9a:	ff_dbi <= 8'h00;
		14'h0a9b:	ff_dbi <= 8'h00;
		14'h0a9c:	ff_dbi <= 8'h00;
		14'h0a9d:	ff_dbi <= 8'h00;
		14'h0a9e:	ff_dbi <= 8'h00;
		14'h0a9f:	ff_dbi <= 8'h00;
		14'h0aa0:	ff_dbi <= 8'h00;
		14'h0aa1:	ff_dbi <= 8'h00;
		14'h0aa2:	ff_dbi <= 8'h00;
		14'h0aa3:	ff_dbi <= 8'h00;
		14'h0aa4:	ff_dbi <= 8'h00;
		14'h0aa5:	ff_dbi <= 8'h00;
		14'h0aa6:	ff_dbi <= 8'h00;
		14'h0aa7:	ff_dbi <= 8'h00;
		14'h0aa8:	ff_dbi <= 8'h00;
		14'h0aa9:	ff_dbi <= 8'h00;
		14'h0aaa:	ff_dbi <= 8'h00;
		14'h0aab:	ff_dbi <= 8'h00;
		14'h0aac:	ff_dbi <= 8'h00;
		14'h0aad:	ff_dbi <= 8'h00;
		14'h0aae:	ff_dbi <= 8'h00;
		14'h0aaf:	ff_dbi <= 8'h00;
		14'h0ab0:	ff_dbi <= 8'h00;
		14'h0ab1:	ff_dbi <= 8'h00;
		14'h0ab2:	ff_dbi <= 8'h00;
		14'h0ab3:	ff_dbi <= 8'h00;
		14'h0ab4:	ff_dbi <= 8'h00;
		14'h0ab5:	ff_dbi <= 8'h00;
		14'h0ab6:	ff_dbi <= 8'h00;
		14'h0ab7:	ff_dbi <= 8'h00;
		14'h0ab8:	ff_dbi <= 8'h00;
		14'h0ab9:	ff_dbi <= 8'h00;
		14'h0aba:	ff_dbi <= 8'h00;
		14'h0abb:	ff_dbi <= 8'h00;
		14'h0abc:	ff_dbi <= 8'h00;
		14'h0abd:	ff_dbi <= 8'h00;
		14'h0abe:	ff_dbi <= 8'h00;
		14'h0abf:	ff_dbi <= 8'h00;
		14'h0ac0:	ff_dbi <= 8'h00;
		14'h0ac1:	ff_dbi <= 8'h00;
		14'h0ac2:	ff_dbi <= 8'h00;
		14'h0ac3:	ff_dbi <= 8'h00;
		14'h0ac4:	ff_dbi <= 8'h00;
		14'h0ac5:	ff_dbi <= 8'h00;
		14'h0ac6:	ff_dbi <= 8'h00;
		14'h0ac7:	ff_dbi <= 8'h00;
		14'h0ac8:	ff_dbi <= 8'h00;
		14'h0ac9:	ff_dbi <= 8'h00;
		14'h0aca:	ff_dbi <= 8'h00;
		14'h0acb:	ff_dbi <= 8'h00;
		14'h0acc:	ff_dbi <= 8'h00;
		14'h0acd:	ff_dbi <= 8'h00;
		14'h0ace:	ff_dbi <= 8'h00;
		14'h0acf:	ff_dbi <= 8'h00;
		14'h0ad0:	ff_dbi <= 8'h00;
		14'h0ad1:	ff_dbi <= 8'h00;
		14'h0ad2:	ff_dbi <= 8'h00;
		14'h0ad3:	ff_dbi <= 8'h00;
		14'h0ad4:	ff_dbi <= 8'h00;
		14'h0ad5:	ff_dbi <= 8'h00;
		14'h0ad6:	ff_dbi <= 8'h00;
		14'h0ad7:	ff_dbi <= 8'h00;
		14'h0ad8:	ff_dbi <= 8'h00;
		14'h0ad9:	ff_dbi <= 8'h00;
		14'h0ada:	ff_dbi <= 8'h00;
		14'h0adb:	ff_dbi <= 8'h00;
		14'h0adc:	ff_dbi <= 8'h00;
		14'h0add:	ff_dbi <= 8'h00;
		14'h0ade:	ff_dbi <= 8'h00;
		14'h0adf:	ff_dbi <= 8'h00;
		14'h0ae0:	ff_dbi <= 8'h00;
		14'h0ae1:	ff_dbi <= 8'h00;
		14'h0ae2:	ff_dbi <= 8'h00;
		14'h0ae3:	ff_dbi <= 8'h00;
		14'h0ae4:	ff_dbi <= 8'h00;
		14'h0ae5:	ff_dbi <= 8'h00;
		14'h0ae6:	ff_dbi <= 8'h00;
		14'h0ae7:	ff_dbi <= 8'h00;
		14'h0ae8:	ff_dbi <= 8'h00;
		14'h0ae9:	ff_dbi <= 8'h00;
		14'h0aea:	ff_dbi <= 8'h00;
		14'h0aeb:	ff_dbi <= 8'h00;
		14'h0aec:	ff_dbi <= 8'h00;
		14'h0aed:	ff_dbi <= 8'h00;
		14'h0aee:	ff_dbi <= 8'h00;
		14'h0aef:	ff_dbi <= 8'h00;
		14'h0af0:	ff_dbi <= 8'h00;
		14'h0af1:	ff_dbi <= 8'h00;
		14'h0af2:	ff_dbi <= 8'h00;
		14'h0af3:	ff_dbi <= 8'h00;
		14'h0af4:	ff_dbi <= 8'h00;
		14'h0af5:	ff_dbi <= 8'h00;
		14'h0af6:	ff_dbi <= 8'h00;
		14'h0af7:	ff_dbi <= 8'h00;
		14'h0af8:	ff_dbi <= 8'h00;
		14'h0af9:	ff_dbi <= 8'h00;
		14'h0afa:	ff_dbi <= 8'h00;
		14'h0afb:	ff_dbi <= 8'h00;
		14'h0afc:	ff_dbi <= 8'h00;
		14'h0afd:	ff_dbi <= 8'h00;
		14'h0afe:	ff_dbi <= 8'h00;
		14'h0aff:	ff_dbi <= 8'h00;
		14'h0b00:	ff_dbi <= 8'h00;
		14'h0b01:	ff_dbi <= 8'h00;
		14'h0b02:	ff_dbi <= 8'h00;
		14'h0b03:	ff_dbi <= 8'h00;
		14'h0b04:	ff_dbi <= 8'h00;
		14'h0b05:	ff_dbi <= 8'h00;
		14'h0b06:	ff_dbi <= 8'h00;
		14'h0b07:	ff_dbi <= 8'h00;
		14'h0b08:	ff_dbi <= 8'h00;
		14'h0b09:	ff_dbi <= 8'h00;
		14'h0b0a:	ff_dbi <= 8'h00;
		14'h0b0b:	ff_dbi <= 8'h00;
		14'h0b0c:	ff_dbi <= 8'h00;
		14'h0b0d:	ff_dbi <= 8'h00;
		14'h0b0e:	ff_dbi <= 8'h00;
		14'h0b0f:	ff_dbi <= 8'h00;
		14'h0b10:	ff_dbi <= 8'h00;
		14'h0b11:	ff_dbi <= 8'h00;
		14'h0b12:	ff_dbi <= 8'h00;
		14'h0b13:	ff_dbi <= 8'h00;
		14'h0b14:	ff_dbi <= 8'h00;
		14'h0b15:	ff_dbi <= 8'h00;
		14'h0b16:	ff_dbi <= 8'h00;
		14'h0b17:	ff_dbi <= 8'h00;
		14'h0b18:	ff_dbi <= 8'h00;
		14'h0b19:	ff_dbi <= 8'h00;
		14'h0b1a:	ff_dbi <= 8'h00;
		14'h0b1b:	ff_dbi <= 8'h00;
		14'h0b1c:	ff_dbi <= 8'h00;
		14'h0b1d:	ff_dbi <= 8'h00;
		14'h0b1e:	ff_dbi <= 8'h00;
		14'h0b1f:	ff_dbi <= 8'h00;
		14'h0b20:	ff_dbi <= 8'h00;
		14'h0b21:	ff_dbi <= 8'h00;
		14'h0b22:	ff_dbi <= 8'h00;
		14'h0b23:	ff_dbi <= 8'h00;
		14'h0b24:	ff_dbi <= 8'h00;
		14'h0b25:	ff_dbi <= 8'h00;
		14'h0b26:	ff_dbi <= 8'h00;
		14'h0b27:	ff_dbi <= 8'h00;
		14'h0b28:	ff_dbi <= 8'h00;
		14'h0b29:	ff_dbi <= 8'h00;
		14'h0b2a:	ff_dbi <= 8'h00;
		14'h0b2b:	ff_dbi <= 8'h00;
		14'h0b2c:	ff_dbi <= 8'h00;
		14'h0b2d:	ff_dbi <= 8'h00;
		14'h0b2e:	ff_dbi <= 8'h00;
		14'h0b2f:	ff_dbi <= 8'h00;
		14'h0b30:	ff_dbi <= 8'h00;
		14'h0b31:	ff_dbi <= 8'h00;
		14'h0b32:	ff_dbi <= 8'h00;
		14'h0b33:	ff_dbi <= 8'h00;
		14'h0b34:	ff_dbi <= 8'h00;
		14'h0b35:	ff_dbi <= 8'h00;
		14'h0b36:	ff_dbi <= 8'h00;
		14'h0b37:	ff_dbi <= 8'h00;
		14'h0b38:	ff_dbi <= 8'h00;
		14'h0b39:	ff_dbi <= 8'h00;
		14'h0b3a:	ff_dbi <= 8'h00;
		14'h0b3b:	ff_dbi <= 8'h00;
		14'h0b3c:	ff_dbi <= 8'h00;
		14'h0b3d:	ff_dbi <= 8'h00;
		14'h0b3e:	ff_dbi <= 8'h00;
		14'h0b3f:	ff_dbi <= 8'h00;
		14'h0b40:	ff_dbi <= 8'h00;
		14'h0b41:	ff_dbi <= 8'h00;
		14'h0b42:	ff_dbi <= 8'h00;
		14'h0b43:	ff_dbi <= 8'h00;
		14'h0b44:	ff_dbi <= 8'h00;
		14'h0b45:	ff_dbi <= 8'h00;
		14'h0b46:	ff_dbi <= 8'h00;
		14'h0b47:	ff_dbi <= 8'h00;
		14'h0b48:	ff_dbi <= 8'h00;
		14'h0b49:	ff_dbi <= 8'h00;
		14'h0b4a:	ff_dbi <= 8'h00;
		14'h0b4b:	ff_dbi <= 8'h00;
		14'h0b4c:	ff_dbi <= 8'h00;
		14'h0b4d:	ff_dbi <= 8'h00;
		14'h0b4e:	ff_dbi <= 8'h00;
		14'h0b4f:	ff_dbi <= 8'h00;
		14'h0b50:	ff_dbi <= 8'h00;
		14'h0b51:	ff_dbi <= 8'h00;
		14'h0b52:	ff_dbi <= 8'h00;
		14'h0b53:	ff_dbi <= 8'h00;
		14'h0b54:	ff_dbi <= 8'h00;
		14'h0b55:	ff_dbi <= 8'h00;
		14'h0b56:	ff_dbi <= 8'h00;
		14'h0b57:	ff_dbi <= 8'h00;
		14'h0b58:	ff_dbi <= 8'h00;
		14'h0b59:	ff_dbi <= 8'h00;
		14'h0b5a:	ff_dbi <= 8'h00;
		14'h0b5b:	ff_dbi <= 8'h00;
		14'h0b5c:	ff_dbi <= 8'h00;
		14'h0b5d:	ff_dbi <= 8'h00;
		14'h0b5e:	ff_dbi <= 8'h00;
		14'h0b5f:	ff_dbi <= 8'h00;
		14'h0b60:	ff_dbi <= 8'h00;
		14'h0b61:	ff_dbi <= 8'h00;
		14'h0b62:	ff_dbi <= 8'h00;
		14'h0b63:	ff_dbi <= 8'h00;
		14'h0b64:	ff_dbi <= 8'h00;
		14'h0b65:	ff_dbi <= 8'h00;
		14'h0b66:	ff_dbi <= 8'h00;
		14'h0b67:	ff_dbi <= 8'h00;
		14'h0b68:	ff_dbi <= 8'h00;
		14'h0b69:	ff_dbi <= 8'h00;
		14'h0b6a:	ff_dbi <= 8'h00;
		14'h0b6b:	ff_dbi <= 8'h00;
		14'h0b6c:	ff_dbi <= 8'h00;
		14'h0b6d:	ff_dbi <= 8'h00;
		14'h0b6e:	ff_dbi <= 8'h00;
		14'h0b6f:	ff_dbi <= 8'h00;
		14'h0b70:	ff_dbi <= 8'h00;
		14'h0b71:	ff_dbi <= 8'h00;
		14'h0b72:	ff_dbi <= 8'h00;
		14'h0b73:	ff_dbi <= 8'h00;
		14'h0b74:	ff_dbi <= 8'h00;
		14'h0b75:	ff_dbi <= 8'h00;
		14'h0b76:	ff_dbi <= 8'h00;
		14'h0b77:	ff_dbi <= 8'h00;
		14'h0b78:	ff_dbi <= 8'h00;
		14'h0b79:	ff_dbi <= 8'h00;
		14'h0b7a:	ff_dbi <= 8'h00;
		14'h0b7b:	ff_dbi <= 8'h00;
		14'h0b7c:	ff_dbi <= 8'h00;
		14'h0b7d:	ff_dbi <= 8'h00;
		14'h0b7e:	ff_dbi <= 8'h00;
		14'h0b7f:	ff_dbi <= 8'h00;
		14'h0b80:	ff_dbi <= 8'h00;
		14'h0b81:	ff_dbi <= 8'h00;
		14'h0b82:	ff_dbi <= 8'h00;
		14'h0b83:	ff_dbi <= 8'h00;
		14'h0b84:	ff_dbi <= 8'h00;
		14'h0b85:	ff_dbi <= 8'h00;
		14'h0b86:	ff_dbi <= 8'h00;
		14'h0b87:	ff_dbi <= 8'h00;
		14'h0b88:	ff_dbi <= 8'h00;
		14'h0b89:	ff_dbi <= 8'h00;
		14'h0b8a:	ff_dbi <= 8'h00;
		14'h0b8b:	ff_dbi <= 8'h00;
		14'h0b8c:	ff_dbi <= 8'h00;
		14'h0b8d:	ff_dbi <= 8'h00;
		14'h0b8e:	ff_dbi <= 8'h00;
		14'h0b8f:	ff_dbi <= 8'h00;
		14'h0b90:	ff_dbi <= 8'h00;
		14'h0b91:	ff_dbi <= 8'h00;
		14'h0b92:	ff_dbi <= 8'h00;
		14'h0b93:	ff_dbi <= 8'h00;
		14'h0b94:	ff_dbi <= 8'h00;
		14'h0b95:	ff_dbi <= 8'h00;
		14'h0b96:	ff_dbi <= 8'h00;
		14'h0b97:	ff_dbi <= 8'h00;
		14'h0b98:	ff_dbi <= 8'h00;
		14'h0b99:	ff_dbi <= 8'h00;
		14'h0b9a:	ff_dbi <= 8'h00;
		14'h0b9b:	ff_dbi <= 8'h00;
		14'h0b9c:	ff_dbi <= 8'h00;
		14'h0b9d:	ff_dbi <= 8'h00;
		14'h0b9e:	ff_dbi <= 8'h00;
		14'h0b9f:	ff_dbi <= 8'h00;
		14'h0ba0:	ff_dbi <= 8'h00;
		14'h0ba1:	ff_dbi <= 8'h00;
		14'h0ba2:	ff_dbi <= 8'h00;
		14'h0ba3:	ff_dbi <= 8'h00;
		14'h0ba4:	ff_dbi <= 8'h00;
		14'h0ba5:	ff_dbi <= 8'h00;
		14'h0ba6:	ff_dbi <= 8'h00;
		14'h0ba7:	ff_dbi <= 8'h00;
		14'h0ba8:	ff_dbi <= 8'h00;
		14'h0ba9:	ff_dbi <= 8'h00;
		14'h0baa:	ff_dbi <= 8'h00;
		14'h0bab:	ff_dbi <= 8'h00;
		14'h0bac:	ff_dbi <= 8'h00;
		14'h0bad:	ff_dbi <= 8'h00;
		14'h0bae:	ff_dbi <= 8'h00;
		14'h0baf:	ff_dbi <= 8'h00;
		14'h0bb0:	ff_dbi <= 8'h00;
		14'h0bb1:	ff_dbi <= 8'h00;
		14'h0bb2:	ff_dbi <= 8'h00;
		14'h0bb3:	ff_dbi <= 8'h00;
		14'h0bb4:	ff_dbi <= 8'h00;
		14'h0bb5:	ff_dbi <= 8'h00;
		14'h0bb6:	ff_dbi <= 8'h00;
		14'h0bb7:	ff_dbi <= 8'h00;
		14'h0bb8:	ff_dbi <= 8'h00;
		14'h0bb9:	ff_dbi <= 8'h00;
		14'h0bba:	ff_dbi <= 8'h00;
		14'h0bbb:	ff_dbi <= 8'h00;
		14'h0bbc:	ff_dbi <= 8'h00;
		14'h0bbd:	ff_dbi <= 8'h00;
		14'h0bbe:	ff_dbi <= 8'h00;
		14'h0bbf:	ff_dbi <= 8'h00;
		14'h0bc0:	ff_dbi <= 8'h00;
		14'h0bc1:	ff_dbi <= 8'h00;
		14'h0bc2:	ff_dbi <= 8'h00;
		14'h0bc3:	ff_dbi <= 8'h00;
		14'h0bc4:	ff_dbi <= 8'h00;
		14'h0bc5:	ff_dbi <= 8'h00;
		14'h0bc6:	ff_dbi <= 8'h00;
		14'h0bc7:	ff_dbi <= 8'h00;
		14'h0bc8:	ff_dbi <= 8'h00;
		14'h0bc9:	ff_dbi <= 8'h00;
		14'h0bca:	ff_dbi <= 8'h00;
		14'h0bcb:	ff_dbi <= 8'h00;
		14'h0bcc:	ff_dbi <= 8'h00;
		14'h0bcd:	ff_dbi <= 8'h00;
		14'h0bce:	ff_dbi <= 8'h00;
		14'h0bcf:	ff_dbi <= 8'h00;
		14'h0bd0:	ff_dbi <= 8'h00;
		14'h0bd1:	ff_dbi <= 8'h00;
		14'h0bd2:	ff_dbi <= 8'h00;
		14'h0bd3:	ff_dbi <= 8'h00;
		14'h0bd4:	ff_dbi <= 8'h00;
		14'h0bd5:	ff_dbi <= 8'h00;
		14'h0bd6:	ff_dbi <= 8'h00;
		14'h0bd7:	ff_dbi <= 8'h00;
		14'h0bd8:	ff_dbi <= 8'h00;
		14'h0bd9:	ff_dbi <= 8'h00;
		14'h0bda:	ff_dbi <= 8'h00;
		14'h0bdb:	ff_dbi <= 8'h00;
		14'h0bdc:	ff_dbi <= 8'h00;
		14'h0bdd:	ff_dbi <= 8'h00;
		14'h0bde:	ff_dbi <= 8'h00;
		14'h0bdf:	ff_dbi <= 8'h00;
		14'h0be0:	ff_dbi <= 8'h00;
		14'h0be1:	ff_dbi <= 8'h00;
		14'h0be2:	ff_dbi <= 8'h00;
		14'h0be3:	ff_dbi <= 8'h00;
		14'h0be4:	ff_dbi <= 8'h00;
		14'h0be5:	ff_dbi <= 8'h00;
		14'h0be6:	ff_dbi <= 8'h00;
		14'h0be7:	ff_dbi <= 8'h00;
		14'h0be8:	ff_dbi <= 8'h00;
		14'h0be9:	ff_dbi <= 8'h00;
		14'h0bea:	ff_dbi <= 8'h00;
		14'h0beb:	ff_dbi <= 8'h00;
		14'h0bec:	ff_dbi <= 8'h00;
		14'h0bed:	ff_dbi <= 8'h00;
		14'h0bee:	ff_dbi <= 8'h00;
		14'h0bef:	ff_dbi <= 8'h00;
		14'h0bf0:	ff_dbi <= 8'h00;
		14'h0bf1:	ff_dbi <= 8'h00;
		14'h0bf2:	ff_dbi <= 8'h00;
		14'h0bf3:	ff_dbi <= 8'h00;
		14'h0bf4:	ff_dbi <= 8'h00;
		14'h0bf5:	ff_dbi <= 8'h00;
		14'h0bf6:	ff_dbi <= 8'h00;
		14'h0bf7:	ff_dbi <= 8'h00;
		14'h0bf8:	ff_dbi <= 8'h00;
		14'h0bf9:	ff_dbi <= 8'h00;
		14'h0bfa:	ff_dbi <= 8'h00;
		14'h0bfb:	ff_dbi <= 8'h00;
		14'h0bfc:	ff_dbi <= 8'h00;
		14'h0bfd:	ff_dbi <= 8'h00;
		14'h0bfe:	ff_dbi <= 8'h00;
		14'h0bff:	ff_dbi <= 8'h00;
		14'h0c00:	ff_dbi <= 8'h00;
		14'h0c01:	ff_dbi <= 8'h00;
		14'h0c02:	ff_dbi <= 8'h00;
		14'h0c03:	ff_dbi <= 8'h00;
		14'h0c04:	ff_dbi <= 8'h00;
		14'h0c05:	ff_dbi <= 8'h00;
		14'h0c06:	ff_dbi <= 8'h00;
		14'h0c07:	ff_dbi <= 8'h00;
		14'h0c08:	ff_dbi <= 8'h00;
		14'h0c09:	ff_dbi <= 8'h00;
		14'h0c0a:	ff_dbi <= 8'h00;
		14'h0c0b:	ff_dbi <= 8'h00;
		14'h0c0c:	ff_dbi <= 8'h00;
		14'h0c0d:	ff_dbi <= 8'h00;
		14'h0c0e:	ff_dbi <= 8'h00;
		14'h0c0f:	ff_dbi <= 8'h00;
		14'h0c10:	ff_dbi <= 8'h00;
		14'h0c11:	ff_dbi <= 8'h00;
		14'h0c12:	ff_dbi <= 8'h00;
		14'h0c13:	ff_dbi <= 8'h00;
		14'h0c14:	ff_dbi <= 8'h00;
		14'h0c15:	ff_dbi <= 8'h00;
		14'h0c16:	ff_dbi <= 8'h00;
		14'h0c17:	ff_dbi <= 8'h00;
		14'h0c18:	ff_dbi <= 8'h00;
		14'h0c19:	ff_dbi <= 8'h00;
		14'h0c1a:	ff_dbi <= 8'h00;
		14'h0c1b:	ff_dbi <= 8'h00;
		14'h0c1c:	ff_dbi <= 8'h00;
		14'h0c1d:	ff_dbi <= 8'h00;
		14'h0c1e:	ff_dbi <= 8'h00;
		14'h0c1f:	ff_dbi <= 8'h00;
		14'h0c20:	ff_dbi <= 8'h00;
		14'h0c21:	ff_dbi <= 8'h00;
		14'h0c22:	ff_dbi <= 8'h00;
		14'h0c23:	ff_dbi <= 8'h00;
		14'h0c24:	ff_dbi <= 8'h00;
		14'h0c25:	ff_dbi <= 8'h00;
		14'h0c26:	ff_dbi <= 8'h00;
		14'h0c27:	ff_dbi <= 8'h00;
		14'h0c28:	ff_dbi <= 8'h00;
		14'h0c29:	ff_dbi <= 8'h00;
		14'h0c2a:	ff_dbi <= 8'h00;
		14'h0c2b:	ff_dbi <= 8'h00;
		14'h0c2c:	ff_dbi <= 8'h00;
		14'h0c2d:	ff_dbi <= 8'h00;
		14'h0c2e:	ff_dbi <= 8'h00;
		14'h0c2f:	ff_dbi <= 8'h00;
		14'h0c30:	ff_dbi <= 8'h00;
		14'h0c31:	ff_dbi <= 8'h00;
		14'h0c32:	ff_dbi <= 8'h00;
		14'h0c33:	ff_dbi <= 8'h00;
		14'h0c34:	ff_dbi <= 8'h00;
		14'h0c35:	ff_dbi <= 8'h00;
		14'h0c36:	ff_dbi <= 8'h00;
		14'h0c37:	ff_dbi <= 8'h00;
		14'h0c38:	ff_dbi <= 8'h00;
		14'h0c39:	ff_dbi <= 8'h00;
		14'h0c3a:	ff_dbi <= 8'h00;
		14'h0c3b:	ff_dbi <= 8'h00;
		14'h0c3c:	ff_dbi <= 8'h00;
		14'h0c3d:	ff_dbi <= 8'h00;
		14'h0c3e:	ff_dbi <= 8'h00;
		14'h0c3f:	ff_dbi <= 8'h00;
		14'h0c40:	ff_dbi <= 8'h00;
		14'h0c41:	ff_dbi <= 8'h00;
		14'h0c42:	ff_dbi <= 8'h00;
		14'h0c43:	ff_dbi <= 8'h00;
		14'h0c44:	ff_dbi <= 8'h00;
		14'h0c45:	ff_dbi <= 8'h00;
		14'h0c46:	ff_dbi <= 8'h00;
		14'h0c47:	ff_dbi <= 8'h00;
		14'h0c48:	ff_dbi <= 8'h00;
		14'h0c49:	ff_dbi <= 8'h00;
		14'h0c4a:	ff_dbi <= 8'h00;
		14'h0c4b:	ff_dbi <= 8'h00;
		14'h0c4c:	ff_dbi <= 8'h00;
		14'h0c4d:	ff_dbi <= 8'h00;
		14'h0c4e:	ff_dbi <= 8'h00;
		14'h0c4f:	ff_dbi <= 8'h00;
		14'h0c50:	ff_dbi <= 8'h00;
		14'h0c51:	ff_dbi <= 8'h00;
		14'h0c52:	ff_dbi <= 8'h00;
		14'h0c53:	ff_dbi <= 8'h00;
		14'h0c54:	ff_dbi <= 8'h00;
		14'h0c55:	ff_dbi <= 8'h00;
		14'h0c56:	ff_dbi <= 8'h00;
		14'h0c57:	ff_dbi <= 8'h00;
		14'h0c58:	ff_dbi <= 8'h00;
		14'h0c59:	ff_dbi <= 8'h00;
		14'h0c5a:	ff_dbi <= 8'h00;
		14'h0c5b:	ff_dbi <= 8'h00;
		14'h0c5c:	ff_dbi <= 8'h00;
		14'h0c5d:	ff_dbi <= 8'h00;
		14'h0c5e:	ff_dbi <= 8'h00;
		14'h0c5f:	ff_dbi <= 8'h00;
		14'h0c60:	ff_dbi <= 8'h00;
		14'h0c61:	ff_dbi <= 8'h00;
		14'h0c62:	ff_dbi <= 8'h00;
		14'h0c63:	ff_dbi <= 8'h00;
		14'h0c64:	ff_dbi <= 8'h00;
		14'h0c65:	ff_dbi <= 8'h00;
		14'h0c66:	ff_dbi <= 8'h00;
		14'h0c67:	ff_dbi <= 8'h00;
		14'h0c68:	ff_dbi <= 8'h00;
		14'h0c69:	ff_dbi <= 8'h00;
		14'h0c6a:	ff_dbi <= 8'h00;
		14'h0c6b:	ff_dbi <= 8'h00;
		14'h0c6c:	ff_dbi <= 8'h00;
		14'h0c6d:	ff_dbi <= 8'h00;
		14'h0c6e:	ff_dbi <= 8'h00;
		14'h0c6f:	ff_dbi <= 8'h00;
		14'h0c70:	ff_dbi <= 8'h00;
		14'h0c71:	ff_dbi <= 8'h00;
		14'h0c72:	ff_dbi <= 8'h00;
		14'h0c73:	ff_dbi <= 8'h00;
		14'h0c74:	ff_dbi <= 8'h00;
		14'h0c75:	ff_dbi <= 8'h00;
		14'h0c76:	ff_dbi <= 8'h00;
		14'h0c77:	ff_dbi <= 8'h00;
		14'h0c78:	ff_dbi <= 8'h00;
		14'h0c79:	ff_dbi <= 8'h00;
		14'h0c7a:	ff_dbi <= 8'h00;
		14'h0c7b:	ff_dbi <= 8'h00;
		14'h0c7c:	ff_dbi <= 8'h00;
		14'h0c7d:	ff_dbi <= 8'h00;
		14'h0c7e:	ff_dbi <= 8'h00;
		14'h0c7f:	ff_dbi <= 8'h00;
		14'h0c80:	ff_dbi <= 8'h00;
		14'h0c81:	ff_dbi <= 8'h00;
		14'h0c82:	ff_dbi <= 8'h00;
		14'h0c83:	ff_dbi <= 8'h00;
		14'h0c84:	ff_dbi <= 8'h00;
		14'h0c85:	ff_dbi <= 8'h00;
		14'h0c86:	ff_dbi <= 8'h00;
		14'h0c87:	ff_dbi <= 8'h00;
		14'h0c88:	ff_dbi <= 8'h00;
		14'h0c89:	ff_dbi <= 8'h00;
		14'h0c8a:	ff_dbi <= 8'h00;
		14'h0c8b:	ff_dbi <= 8'h00;
		14'h0c8c:	ff_dbi <= 8'h00;
		14'h0c8d:	ff_dbi <= 8'h00;
		14'h0c8e:	ff_dbi <= 8'h00;
		14'h0c8f:	ff_dbi <= 8'h00;
		14'h0c90:	ff_dbi <= 8'h00;
		14'h0c91:	ff_dbi <= 8'h00;
		14'h0c92:	ff_dbi <= 8'h00;
		14'h0c93:	ff_dbi <= 8'h00;
		14'h0c94:	ff_dbi <= 8'h00;
		14'h0c95:	ff_dbi <= 8'h00;
		14'h0c96:	ff_dbi <= 8'h00;
		14'h0c97:	ff_dbi <= 8'h00;
		14'h0c98:	ff_dbi <= 8'h00;
		14'h0c99:	ff_dbi <= 8'h00;
		14'h0c9a:	ff_dbi <= 8'h00;
		14'h0c9b:	ff_dbi <= 8'h00;
		14'h0c9c:	ff_dbi <= 8'h00;
		14'h0c9d:	ff_dbi <= 8'h00;
		14'h0c9e:	ff_dbi <= 8'h00;
		14'h0c9f:	ff_dbi <= 8'h00;
		14'h0ca0:	ff_dbi <= 8'h00;
		14'h0ca1:	ff_dbi <= 8'h00;
		14'h0ca2:	ff_dbi <= 8'h00;
		14'h0ca3:	ff_dbi <= 8'h00;
		14'h0ca4:	ff_dbi <= 8'h00;
		14'h0ca5:	ff_dbi <= 8'h00;
		14'h0ca6:	ff_dbi <= 8'h00;
		14'h0ca7:	ff_dbi <= 8'h00;
		14'h0ca8:	ff_dbi <= 8'h00;
		14'h0ca9:	ff_dbi <= 8'h00;
		14'h0caa:	ff_dbi <= 8'h00;
		14'h0cab:	ff_dbi <= 8'h00;
		14'h0cac:	ff_dbi <= 8'h00;
		14'h0cad:	ff_dbi <= 8'h00;
		14'h0cae:	ff_dbi <= 8'h00;
		14'h0caf:	ff_dbi <= 8'h00;
		14'h0cb0:	ff_dbi <= 8'h00;
		14'h0cb1:	ff_dbi <= 8'h00;
		14'h0cb2:	ff_dbi <= 8'h00;
		14'h0cb3:	ff_dbi <= 8'h00;
		14'h0cb4:	ff_dbi <= 8'h00;
		14'h0cb5:	ff_dbi <= 8'h00;
		14'h0cb6:	ff_dbi <= 8'h00;
		14'h0cb7:	ff_dbi <= 8'h00;
		14'h0cb8:	ff_dbi <= 8'h00;
		14'h0cb9:	ff_dbi <= 8'h00;
		14'h0cba:	ff_dbi <= 8'h00;
		14'h0cbb:	ff_dbi <= 8'h00;
		14'h0cbc:	ff_dbi <= 8'h00;
		14'h0cbd:	ff_dbi <= 8'h00;
		14'h0cbe:	ff_dbi <= 8'h00;
		14'h0cbf:	ff_dbi <= 8'h00;
		14'h0cc0:	ff_dbi <= 8'h00;
		14'h0cc1:	ff_dbi <= 8'h00;
		14'h0cc2:	ff_dbi <= 8'h00;
		14'h0cc3:	ff_dbi <= 8'h00;
		14'h0cc4:	ff_dbi <= 8'h00;
		14'h0cc5:	ff_dbi <= 8'h00;
		14'h0cc6:	ff_dbi <= 8'h00;
		14'h0cc7:	ff_dbi <= 8'h00;
		14'h0cc8:	ff_dbi <= 8'h00;
		14'h0cc9:	ff_dbi <= 8'h00;
		14'h0cca:	ff_dbi <= 8'h00;
		14'h0ccb:	ff_dbi <= 8'h00;
		14'h0ccc:	ff_dbi <= 8'h00;
		14'h0ccd:	ff_dbi <= 8'h00;
		14'h0cce:	ff_dbi <= 8'h00;
		14'h0ccf:	ff_dbi <= 8'h00;
		14'h0cd0:	ff_dbi <= 8'h00;
		14'h0cd1:	ff_dbi <= 8'h00;
		14'h0cd2:	ff_dbi <= 8'h00;
		14'h0cd3:	ff_dbi <= 8'h00;
		14'h0cd4:	ff_dbi <= 8'h00;
		14'h0cd5:	ff_dbi <= 8'h00;
		14'h0cd6:	ff_dbi <= 8'h00;
		14'h0cd7:	ff_dbi <= 8'h00;
		14'h0cd8:	ff_dbi <= 8'h00;
		14'h0cd9:	ff_dbi <= 8'h00;
		14'h0cda:	ff_dbi <= 8'h00;
		14'h0cdb:	ff_dbi <= 8'h00;
		14'h0cdc:	ff_dbi <= 8'h00;
		14'h0cdd:	ff_dbi <= 8'h00;
		14'h0cde:	ff_dbi <= 8'h00;
		14'h0cdf:	ff_dbi <= 8'h00;
		14'h0ce0:	ff_dbi <= 8'h00;
		14'h0ce1:	ff_dbi <= 8'h00;
		14'h0ce2:	ff_dbi <= 8'h00;
		14'h0ce3:	ff_dbi <= 8'h00;
		14'h0ce4:	ff_dbi <= 8'h00;
		14'h0ce5:	ff_dbi <= 8'h00;
		14'h0ce6:	ff_dbi <= 8'h00;
		14'h0ce7:	ff_dbi <= 8'h00;
		14'h0ce8:	ff_dbi <= 8'h00;
		14'h0ce9:	ff_dbi <= 8'h00;
		14'h0cea:	ff_dbi <= 8'h00;
		14'h0ceb:	ff_dbi <= 8'h00;
		14'h0cec:	ff_dbi <= 8'h00;
		14'h0ced:	ff_dbi <= 8'h00;
		14'h0cee:	ff_dbi <= 8'h00;
		14'h0cef:	ff_dbi <= 8'h00;
		14'h0cf0:	ff_dbi <= 8'h00;
		14'h0cf1:	ff_dbi <= 8'h00;
		14'h0cf2:	ff_dbi <= 8'h00;
		14'h0cf3:	ff_dbi <= 8'h00;
		14'h0cf4:	ff_dbi <= 8'h00;
		14'h0cf5:	ff_dbi <= 8'h00;
		14'h0cf6:	ff_dbi <= 8'h00;
		14'h0cf7:	ff_dbi <= 8'h00;
		14'h0cf8:	ff_dbi <= 8'h00;
		14'h0cf9:	ff_dbi <= 8'h00;
		14'h0cfa:	ff_dbi <= 8'h00;
		14'h0cfb:	ff_dbi <= 8'h00;
		14'h0cfc:	ff_dbi <= 8'h00;
		14'h0cfd:	ff_dbi <= 8'h00;
		14'h0cfe:	ff_dbi <= 8'h00;
		14'h0cff:	ff_dbi <= 8'h00;
		14'h0d00:	ff_dbi <= 8'h00;
		14'h0d01:	ff_dbi <= 8'h00;
		14'h0d02:	ff_dbi <= 8'h00;
		14'h0d03:	ff_dbi <= 8'h00;
		14'h0d04:	ff_dbi <= 8'h00;
		14'h0d05:	ff_dbi <= 8'h00;
		14'h0d06:	ff_dbi <= 8'h00;
		14'h0d07:	ff_dbi <= 8'h00;
		14'h0d08:	ff_dbi <= 8'h00;
		14'h0d09:	ff_dbi <= 8'h00;
		14'h0d0a:	ff_dbi <= 8'h00;
		14'h0d0b:	ff_dbi <= 8'h00;
		14'h0d0c:	ff_dbi <= 8'h00;
		14'h0d0d:	ff_dbi <= 8'h00;
		14'h0d0e:	ff_dbi <= 8'h00;
		14'h0d0f:	ff_dbi <= 8'h00;
		14'h0d10:	ff_dbi <= 8'h00;
		14'h0d11:	ff_dbi <= 8'h00;
		14'h0d12:	ff_dbi <= 8'h00;
		14'h0d13:	ff_dbi <= 8'h00;
		14'h0d14:	ff_dbi <= 8'h00;
		14'h0d15:	ff_dbi <= 8'h00;
		14'h0d16:	ff_dbi <= 8'h00;
		14'h0d17:	ff_dbi <= 8'h00;
		14'h0d18:	ff_dbi <= 8'h00;
		14'h0d19:	ff_dbi <= 8'h00;
		14'h0d1a:	ff_dbi <= 8'h00;
		14'h0d1b:	ff_dbi <= 8'h00;
		14'h0d1c:	ff_dbi <= 8'h00;
		14'h0d1d:	ff_dbi <= 8'h00;
		14'h0d1e:	ff_dbi <= 8'h00;
		14'h0d1f:	ff_dbi <= 8'h00;
		14'h0d20:	ff_dbi <= 8'h00;
		14'h0d21:	ff_dbi <= 8'h00;
		14'h0d22:	ff_dbi <= 8'h00;
		14'h0d23:	ff_dbi <= 8'h00;
		14'h0d24:	ff_dbi <= 8'h00;
		14'h0d25:	ff_dbi <= 8'h00;
		14'h0d26:	ff_dbi <= 8'h00;
		14'h0d27:	ff_dbi <= 8'h00;
		14'h0d28:	ff_dbi <= 8'h00;
		14'h0d29:	ff_dbi <= 8'h00;
		14'h0d2a:	ff_dbi <= 8'h00;
		14'h0d2b:	ff_dbi <= 8'h00;
		14'h0d2c:	ff_dbi <= 8'h00;
		14'h0d2d:	ff_dbi <= 8'h00;
		14'h0d2e:	ff_dbi <= 8'h00;
		14'h0d2f:	ff_dbi <= 8'h00;
		14'h0d30:	ff_dbi <= 8'h00;
		14'h0d31:	ff_dbi <= 8'h00;
		14'h0d32:	ff_dbi <= 8'h00;
		14'h0d33:	ff_dbi <= 8'h00;
		14'h0d34:	ff_dbi <= 8'h00;
		14'h0d35:	ff_dbi <= 8'h00;
		14'h0d36:	ff_dbi <= 8'h00;
		14'h0d37:	ff_dbi <= 8'h00;
		14'h0d38:	ff_dbi <= 8'h00;
		14'h0d39:	ff_dbi <= 8'h00;
		14'h0d3a:	ff_dbi <= 8'h00;
		14'h0d3b:	ff_dbi <= 8'h00;
		14'h0d3c:	ff_dbi <= 8'h00;
		14'h0d3d:	ff_dbi <= 8'h00;
		14'h0d3e:	ff_dbi <= 8'h00;
		14'h0d3f:	ff_dbi <= 8'h00;
		14'h0d40:	ff_dbi <= 8'h00;
		14'h0d41:	ff_dbi <= 8'h00;
		14'h0d42:	ff_dbi <= 8'h00;
		14'h0d43:	ff_dbi <= 8'h00;
		14'h0d44:	ff_dbi <= 8'h00;
		14'h0d45:	ff_dbi <= 8'h00;
		14'h0d46:	ff_dbi <= 8'h00;
		14'h0d47:	ff_dbi <= 8'h00;
		14'h0d48:	ff_dbi <= 8'h00;
		14'h0d49:	ff_dbi <= 8'h00;
		14'h0d4a:	ff_dbi <= 8'h00;
		14'h0d4b:	ff_dbi <= 8'h00;
		14'h0d4c:	ff_dbi <= 8'h00;
		14'h0d4d:	ff_dbi <= 8'h00;
		14'h0d4e:	ff_dbi <= 8'h00;
		14'h0d4f:	ff_dbi <= 8'h00;
		14'h0d50:	ff_dbi <= 8'h00;
		14'h0d51:	ff_dbi <= 8'h00;
		14'h0d52:	ff_dbi <= 8'h00;
		14'h0d53:	ff_dbi <= 8'h00;
		14'h0d54:	ff_dbi <= 8'h00;
		14'h0d55:	ff_dbi <= 8'h00;
		14'h0d56:	ff_dbi <= 8'h00;
		14'h0d57:	ff_dbi <= 8'h00;
		14'h0d58:	ff_dbi <= 8'h00;
		14'h0d59:	ff_dbi <= 8'h00;
		14'h0d5a:	ff_dbi <= 8'h00;
		14'h0d5b:	ff_dbi <= 8'h00;
		14'h0d5c:	ff_dbi <= 8'h00;
		14'h0d5d:	ff_dbi <= 8'h00;
		14'h0d5e:	ff_dbi <= 8'h00;
		14'h0d5f:	ff_dbi <= 8'h00;
		14'h0d60:	ff_dbi <= 8'h00;
		14'h0d61:	ff_dbi <= 8'h00;
		14'h0d62:	ff_dbi <= 8'h00;
		14'h0d63:	ff_dbi <= 8'h00;
		14'h0d64:	ff_dbi <= 8'h00;
		14'h0d65:	ff_dbi <= 8'h00;
		14'h0d66:	ff_dbi <= 8'h00;
		14'h0d67:	ff_dbi <= 8'h00;
		14'h0d68:	ff_dbi <= 8'h00;
		14'h0d69:	ff_dbi <= 8'h00;
		14'h0d6a:	ff_dbi <= 8'h00;
		14'h0d6b:	ff_dbi <= 8'h00;
		14'h0d6c:	ff_dbi <= 8'h00;
		14'h0d6d:	ff_dbi <= 8'h00;
		14'h0d6e:	ff_dbi <= 8'h00;
		14'h0d6f:	ff_dbi <= 8'h00;
		14'h0d70:	ff_dbi <= 8'h00;
		14'h0d71:	ff_dbi <= 8'h00;
		14'h0d72:	ff_dbi <= 8'h00;
		14'h0d73:	ff_dbi <= 8'h00;
		14'h0d74:	ff_dbi <= 8'h00;
		14'h0d75:	ff_dbi <= 8'h00;
		14'h0d76:	ff_dbi <= 8'h00;
		14'h0d77:	ff_dbi <= 8'h00;
		14'h0d78:	ff_dbi <= 8'h00;
		14'h0d79:	ff_dbi <= 8'h00;
		14'h0d7a:	ff_dbi <= 8'h00;
		14'h0d7b:	ff_dbi <= 8'h00;
		14'h0d7c:	ff_dbi <= 8'h00;
		14'h0d7d:	ff_dbi <= 8'h00;
		14'h0d7e:	ff_dbi <= 8'h00;
		14'h0d7f:	ff_dbi <= 8'h00;
		14'h0d80:	ff_dbi <= 8'h00;
		14'h0d81:	ff_dbi <= 8'h00;
		14'h0d82:	ff_dbi <= 8'h00;
		14'h0d83:	ff_dbi <= 8'h00;
		14'h0d84:	ff_dbi <= 8'h00;
		14'h0d85:	ff_dbi <= 8'h00;
		14'h0d86:	ff_dbi <= 8'h00;
		14'h0d87:	ff_dbi <= 8'h00;
		14'h0d88:	ff_dbi <= 8'h00;
		14'h0d89:	ff_dbi <= 8'h00;
		14'h0d8a:	ff_dbi <= 8'h00;
		14'h0d8b:	ff_dbi <= 8'h00;
		14'h0d8c:	ff_dbi <= 8'h00;
		14'h0d8d:	ff_dbi <= 8'h00;
		14'h0d8e:	ff_dbi <= 8'h00;
		14'h0d8f:	ff_dbi <= 8'h00;
		14'h0d90:	ff_dbi <= 8'h00;
		14'h0d91:	ff_dbi <= 8'h00;
		14'h0d92:	ff_dbi <= 8'h00;
		14'h0d93:	ff_dbi <= 8'h00;
		14'h0d94:	ff_dbi <= 8'h00;
		14'h0d95:	ff_dbi <= 8'h00;
		14'h0d96:	ff_dbi <= 8'h00;
		14'h0d97:	ff_dbi <= 8'h00;
		14'h0d98:	ff_dbi <= 8'h00;
		14'h0d99:	ff_dbi <= 8'h00;
		14'h0d9a:	ff_dbi <= 8'h00;
		14'h0d9b:	ff_dbi <= 8'h00;
		14'h0d9c:	ff_dbi <= 8'h00;
		14'h0d9d:	ff_dbi <= 8'h00;
		14'h0d9e:	ff_dbi <= 8'h00;
		14'h0d9f:	ff_dbi <= 8'h00;
		14'h0da0:	ff_dbi <= 8'h00;
		14'h0da1:	ff_dbi <= 8'h00;
		14'h0da2:	ff_dbi <= 8'h00;
		14'h0da3:	ff_dbi <= 8'h00;
		14'h0da4:	ff_dbi <= 8'h00;
		14'h0da5:	ff_dbi <= 8'h00;
		14'h0da6:	ff_dbi <= 8'h00;
		14'h0da7:	ff_dbi <= 8'h00;
		14'h0da8:	ff_dbi <= 8'h00;
		14'h0da9:	ff_dbi <= 8'h00;
		14'h0daa:	ff_dbi <= 8'h00;
		14'h0dab:	ff_dbi <= 8'h00;
		14'h0dac:	ff_dbi <= 8'h00;
		14'h0dad:	ff_dbi <= 8'h00;
		14'h0dae:	ff_dbi <= 8'h00;
		14'h0daf:	ff_dbi <= 8'h00;
		14'h0db0:	ff_dbi <= 8'h00;
		14'h0db1:	ff_dbi <= 8'h00;
		14'h0db2:	ff_dbi <= 8'h00;
		14'h0db3:	ff_dbi <= 8'h00;
		14'h0db4:	ff_dbi <= 8'h00;
		14'h0db5:	ff_dbi <= 8'h00;
		14'h0db6:	ff_dbi <= 8'h00;
		14'h0db7:	ff_dbi <= 8'h00;
		14'h0db8:	ff_dbi <= 8'h00;
		14'h0db9:	ff_dbi <= 8'h00;
		14'h0dba:	ff_dbi <= 8'h00;
		14'h0dbb:	ff_dbi <= 8'h00;
		14'h0dbc:	ff_dbi <= 8'h00;
		14'h0dbd:	ff_dbi <= 8'h00;
		14'h0dbe:	ff_dbi <= 8'h00;
		14'h0dbf:	ff_dbi <= 8'h00;
		14'h0dc0:	ff_dbi <= 8'h00;
		14'h0dc1:	ff_dbi <= 8'h00;
		14'h0dc2:	ff_dbi <= 8'h00;
		14'h0dc3:	ff_dbi <= 8'h00;
		14'h0dc4:	ff_dbi <= 8'h00;
		14'h0dc5:	ff_dbi <= 8'h00;
		14'h0dc6:	ff_dbi <= 8'h00;
		14'h0dc7:	ff_dbi <= 8'h00;
		14'h0dc8:	ff_dbi <= 8'h00;
		14'h0dc9:	ff_dbi <= 8'h00;
		14'h0dca:	ff_dbi <= 8'h00;
		14'h0dcb:	ff_dbi <= 8'h00;
		14'h0dcc:	ff_dbi <= 8'h00;
		14'h0dcd:	ff_dbi <= 8'h00;
		14'h0dce:	ff_dbi <= 8'h00;
		14'h0dcf:	ff_dbi <= 8'h00;
		14'h0dd0:	ff_dbi <= 8'h00;
		14'h0dd1:	ff_dbi <= 8'h00;
		14'h0dd2:	ff_dbi <= 8'h00;
		14'h0dd3:	ff_dbi <= 8'h00;
		14'h0dd4:	ff_dbi <= 8'h00;
		14'h0dd5:	ff_dbi <= 8'h00;
		14'h0dd6:	ff_dbi <= 8'h00;
		14'h0dd7:	ff_dbi <= 8'h00;
		14'h0dd8:	ff_dbi <= 8'h00;
		14'h0dd9:	ff_dbi <= 8'h00;
		14'h0dda:	ff_dbi <= 8'h00;
		14'h0ddb:	ff_dbi <= 8'h00;
		14'h0ddc:	ff_dbi <= 8'h00;
		14'h0ddd:	ff_dbi <= 8'h00;
		14'h0dde:	ff_dbi <= 8'h00;
		14'h0ddf:	ff_dbi <= 8'h00;
		14'h0de0:	ff_dbi <= 8'h00;
		14'h0de1:	ff_dbi <= 8'h00;
		14'h0de2:	ff_dbi <= 8'h00;
		14'h0de3:	ff_dbi <= 8'h00;
		14'h0de4:	ff_dbi <= 8'h00;
		14'h0de5:	ff_dbi <= 8'h00;
		14'h0de6:	ff_dbi <= 8'h00;
		14'h0de7:	ff_dbi <= 8'h00;
		14'h0de8:	ff_dbi <= 8'h00;
		14'h0de9:	ff_dbi <= 8'h00;
		14'h0dea:	ff_dbi <= 8'h00;
		14'h0deb:	ff_dbi <= 8'h00;
		14'h0dec:	ff_dbi <= 8'h00;
		14'h0ded:	ff_dbi <= 8'h00;
		14'h0dee:	ff_dbi <= 8'h00;
		14'h0def:	ff_dbi <= 8'h00;
		14'h0df0:	ff_dbi <= 8'h00;
		14'h0df1:	ff_dbi <= 8'h00;
		14'h0df2:	ff_dbi <= 8'h00;
		14'h0df3:	ff_dbi <= 8'h00;
		14'h0df4:	ff_dbi <= 8'h00;
		14'h0df5:	ff_dbi <= 8'h00;
		14'h0df6:	ff_dbi <= 8'h00;
		14'h0df7:	ff_dbi <= 8'h00;
		14'h0df8:	ff_dbi <= 8'h00;
		14'h0df9:	ff_dbi <= 8'h00;
		14'h0dfa:	ff_dbi <= 8'h00;
		14'h0dfb:	ff_dbi <= 8'h00;
		14'h0dfc:	ff_dbi <= 8'h00;
		14'h0dfd:	ff_dbi <= 8'h00;
		14'h0dfe:	ff_dbi <= 8'h00;
		14'h0dff:	ff_dbi <= 8'h00;
		14'h0e00:	ff_dbi <= 8'h00;
		14'h0e01:	ff_dbi <= 8'h00;
		14'h0e02:	ff_dbi <= 8'h00;
		14'h0e03:	ff_dbi <= 8'h00;
		14'h0e04:	ff_dbi <= 8'h00;
		14'h0e05:	ff_dbi <= 8'h00;
		14'h0e06:	ff_dbi <= 8'h00;
		14'h0e07:	ff_dbi <= 8'h00;
		14'h0e08:	ff_dbi <= 8'h00;
		14'h0e09:	ff_dbi <= 8'h00;
		14'h0e0a:	ff_dbi <= 8'h00;
		14'h0e0b:	ff_dbi <= 8'h00;
		14'h0e0c:	ff_dbi <= 8'h00;
		14'h0e0d:	ff_dbi <= 8'h00;
		14'h0e0e:	ff_dbi <= 8'h00;
		14'h0e0f:	ff_dbi <= 8'h00;
		14'h0e10:	ff_dbi <= 8'h00;
		14'h0e11:	ff_dbi <= 8'h00;
		14'h0e12:	ff_dbi <= 8'h00;
		14'h0e13:	ff_dbi <= 8'h00;
		14'h0e14:	ff_dbi <= 8'h00;
		14'h0e15:	ff_dbi <= 8'h00;
		14'h0e16:	ff_dbi <= 8'h00;
		14'h0e17:	ff_dbi <= 8'h00;
		14'h0e18:	ff_dbi <= 8'h00;
		14'h0e19:	ff_dbi <= 8'h00;
		14'h0e1a:	ff_dbi <= 8'h00;
		14'h0e1b:	ff_dbi <= 8'h00;
		14'h0e1c:	ff_dbi <= 8'h00;
		14'h0e1d:	ff_dbi <= 8'h00;
		14'h0e1e:	ff_dbi <= 8'h00;
		14'h0e1f:	ff_dbi <= 8'h00;
		14'h0e20:	ff_dbi <= 8'h00;
		14'h0e21:	ff_dbi <= 8'h00;
		14'h0e22:	ff_dbi <= 8'h00;
		14'h0e23:	ff_dbi <= 8'h00;
		14'h0e24:	ff_dbi <= 8'h00;
		14'h0e25:	ff_dbi <= 8'h00;
		14'h0e26:	ff_dbi <= 8'h00;
		14'h0e27:	ff_dbi <= 8'h00;
		14'h0e28:	ff_dbi <= 8'h00;
		14'h0e29:	ff_dbi <= 8'h00;
		14'h0e2a:	ff_dbi <= 8'h00;
		14'h0e2b:	ff_dbi <= 8'h00;
		14'h0e2c:	ff_dbi <= 8'h00;
		14'h0e2d:	ff_dbi <= 8'h00;
		14'h0e2e:	ff_dbi <= 8'h00;
		14'h0e2f:	ff_dbi <= 8'h00;
		14'h0e30:	ff_dbi <= 8'h00;
		14'h0e31:	ff_dbi <= 8'h00;
		14'h0e32:	ff_dbi <= 8'h00;
		14'h0e33:	ff_dbi <= 8'h00;
		14'h0e34:	ff_dbi <= 8'h00;
		14'h0e35:	ff_dbi <= 8'h00;
		14'h0e36:	ff_dbi <= 8'h00;
		14'h0e37:	ff_dbi <= 8'h00;
		14'h0e38:	ff_dbi <= 8'h00;
		14'h0e39:	ff_dbi <= 8'h00;
		14'h0e3a:	ff_dbi <= 8'h00;
		14'h0e3b:	ff_dbi <= 8'h00;
		14'h0e3c:	ff_dbi <= 8'h00;
		14'h0e3d:	ff_dbi <= 8'h00;
		14'h0e3e:	ff_dbi <= 8'h00;
		14'h0e3f:	ff_dbi <= 8'h00;
		14'h0e40:	ff_dbi <= 8'h00;
		14'h0e41:	ff_dbi <= 8'h00;
		14'h0e42:	ff_dbi <= 8'h00;
		14'h0e43:	ff_dbi <= 8'h00;
		14'h0e44:	ff_dbi <= 8'h00;
		14'h0e45:	ff_dbi <= 8'h00;
		14'h0e46:	ff_dbi <= 8'h00;
		14'h0e47:	ff_dbi <= 8'h00;
		14'h0e48:	ff_dbi <= 8'h00;
		14'h0e49:	ff_dbi <= 8'h00;
		14'h0e4a:	ff_dbi <= 8'h00;
		14'h0e4b:	ff_dbi <= 8'h00;
		14'h0e4c:	ff_dbi <= 8'h00;
		14'h0e4d:	ff_dbi <= 8'h00;
		14'h0e4e:	ff_dbi <= 8'h00;
		14'h0e4f:	ff_dbi <= 8'h00;
		14'h0e50:	ff_dbi <= 8'h00;
		14'h0e51:	ff_dbi <= 8'h00;
		14'h0e52:	ff_dbi <= 8'h00;
		14'h0e53:	ff_dbi <= 8'h00;
		14'h0e54:	ff_dbi <= 8'h00;
		14'h0e55:	ff_dbi <= 8'h00;
		14'h0e56:	ff_dbi <= 8'h00;
		14'h0e57:	ff_dbi <= 8'h00;
		14'h0e58:	ff_dbi <= 8'h00;
		14'h0e59:	ff_dbi <= 8'h00;
		14'h0e5a:	ff_dbi <= 8'h00;
		14'h0e5b:	ff_dbi <= 8'h00;
		14'h0e5c:	ff_dbi <= 8'h00;
		14'h0e5d:	ff_dbi <= 8'h00;
		14'h0e5e:	ff_dbi <= 8'h00;
		14'h0e5f:	ff_dbi <= 8'h00;
		14'h0e60:	ff_dbi <= 8'h00;
		14'h0e61:	ff_dbi <= 8'h00;
		14'h0e62:	ff_dbi <= 8'h00;
		14'h0e63:	ff_dbi <= 8'h00;
		14'h0e64:	ff_dbi <= 8'h00;
		14'h0e65:	ff_dbi <= 8'h00;
		14'h0e66:	ff_dbi <= 8'h00;
		14'h0e67:	ff_dbi <= 8'h00;
		14'h0e68:	ff_dbi <= 8'h00;
		14'h0e69:	ff_dbi <= 8'h00;
		14'h0e6a:	ff_dbi <= 8'h00;
		14'h0e6b:	ff_dbi <= 8'h00;
		14'h0e6c:	ff_dbi <= 8'h00;
		14'h0e6d:	ff_dbi <= 8'h00;
		14'h0e6e:	ff_dbi <= 8'h00;
		14'h0e6f:	ff_dbi <= 8'h00;
		14'h0e70:	ff_dbi <= 8'h00;
		14'h0e71:	ff_dbi <= 8'h00;
		14'h0e72:	ff_dbi <= 8'h00;
		14'h0e73:	ff_dbi <= 8'h00;
		14'h0e74:	ff_dbi <= 8'h00;
		14'h0e75:	ff_dbi <= 8'h00;
		14'h0e76:	ff_dbi <= 8'h00;
		14'h0e77:	ff_dbi <= 8'h00;
		14'h0e78:	ff_dbi <= 8'h00;
		14'h0e79:	ff_dbi <= 8'h00;
		14'h0e7a:	ff_dbi <= 8'h00;
		14'h0e7b:	ff_dbi <= 8'h00;
		14'h0e7c:	ff_dbi <= 8'h00;
		14'h0e7d:	ff_dbi <= 8'h00;
		14'h0e7e:	ff_dbi <= 8'h00;
		14'h0e7f:	ff_dbi <= 8'h00;
		14'h0e80:	ff_dbi <= 8'h00;
		14'h0e81:	ff_dbi <= 8'h00;
		14'h0e82:	ff_dbi <= 8'h00;
		14'h0e83:	ff_dbi <= 8'h00;
		14'h0e84:	ff_dbi <= 8'h00;
		14'h0e85:	ff_dbi <= 8'h00;
		14'h0e86:	ff_dbi <= 8'h00;
		14'h0e87:	ff_dbi <= 8'h00;
		14'h0e88:	ff_dbi <= 8'h00;
		14'h0e89:	ff_dbi <= 8'h00;
		14'h0e8a:	ff_dbi <= 8'h00;
		14'h0e8b:	ff_dbi <= 8'h00;
		14'h0e8c:	ff_dbi <= 8'h00;
		14'h0e8d:	ff_dbi <= 8'h00;
		14'h0e8e:	ff_dbi <= 8'h00;
		14'h0e8f:	ff_dbi <= 8'h00;
		14'h0e90:	ff_dbi <= 8'h00;
		14'h0e91:	ff_dbi <= 8'h00;
		14'h0e92:	ff_dbi <= 8'h00;
		14'h0e93:	ff_dbi <= 8'h00;
		14'h0e94:	ff_dbi <= 8'h00;
		14'h0e95:	ff_dbi <= 8'h00;
		14'h0e96:	ff_dbi <= 8'h00;
		14'h0e97:	ff_dbi <= 8'h00;
		14'h0e98:	ff_dbi <= 8'h00;
		14'h0e99:	ff_dbi <= 8'h00;
		14'h0e9a:	ff_dbi <= 8'h00;
		14'h0e9b:	ff_dbi <= 8'h00;
		14'h0e9c:	ff_dbi <= 8'h00;
		14'h0e9d:	ff_dbi <= 8'h00;
		14'h0e9e:	ff_dbi <= 8'h00;
		14'h0e9f:	ff_dbi <= 8'h00;
		14'h0ea0:	ff_dbi <= 8'h00;
		14'h0ea1:	ff_dbi <= 8'h00;
		14'h0ea2:	ff_dbi <= 8'h00;
		14'h0ea3:	ff_dbi <= 8'h00;
		14'h0ea4:	ff_dbi <= 8'h00;
		14'h0ea5:	ff_dbi <= 8'h00;
		14'h0ea6:	ff_dbi <= 8'h00;
		14'h0ea7:	ff_dbi <= 8'h00;
		14'h0ea8:	ff_dbi <= 8'h00;
		14'h0ea9:	ff_dbi <= 8'h00;
		14'h0eaa:	ff_dbi <= 8'h00;
		14'h0eab:	ff_dbi <= 8'h00;
		14'h0eac:	ff_dbi <= 8'h00;
		14'h0ead:	ff_dbi <= 8'h00;
		14'h0eae:	ff_dbi <= 8'h00;
		14'h0eaf:	ff_dbi <= 8'h00;
		14'h0eb0:	ff_dbi <= 8'h00;
		14'h0eb1:	ff_dbi <= 8'h00;
		14'h0eb2:	ff_dbi <= 8'h00;
		14'h0eb3:	ff_dbi <= 8'h00;
		14'h0eb4:	ff_dbi <= 8'h00;
		14'h0eb5:	ff_dbi <= 8'h00;
		14'h0eb6:	ff_dbi <= 8'h00;
		14'h0eb7:	ff_dbi <= 8'h00;
		14'h0eb8:	ff_dbi <= 8'h00;
		14'h0eb9:	ff_dbi <= 8'h00;
		14'h0eba:	ff_dbi <= 8'h00;
		14'h0ebb:	ff_dbi <= 8'h00;
		14'h0ebc:	ff_dbi <= 8'h00;
		14'h0ebd:	ff_dbi <= 8'h00;
		14'h0ebe:	ff_dbi <= 8'h00;
		14'h0ebf:	ff_dbi <= 8'h00;
		14'h0ec0:	ff_dbi <= 8'h00;
		14'h0ec1:	ff_dbi <= 8'h00;
		14'h0ec2:	ff_dbi <= 8'h00;
		14'h0ec3:	ff_dbi <= 8'h00;
		14'h0ec4:	ff_dbi <= 8'h00;
		14'h0ec5:	ff_dbi <= 8'h00;
		14'h0ec6:	ff_dbi <= 8'h00;
		14'h0ec7:	ff_dbi <= 8'h00;
		14'h0ec8:	ff_dbi <= 8'h00;
		14'h0ec9:	ff_dbi <= 8'h00;
		14'h0eca:	ff_dbi <= 8'h00;
		14'h0ecb:	ff_dbi <= 8'h00;
		14'h0ecc:	ff_dbi <= 8'h00;
		14'h0ecd:	ff_dbi <= 8'h00;
		14'h0ece:	ff_dbi <= 8'h00;
		14'h0ecf:	ff_dbi <= 8'h00;
		14'h0ed0:	ff_dbi <= 8'h00;
		14'h0ed1:	ff_dbi <= 8'h00;
		14'h0ed2:	ff_dbi <= 8'h00;
		14'h0ed3:	ff_dbi <= 8'h00;
		14'h0ed4:	ff_dbi <= 8'h00;
		14'h0ed5:	ff_dbi <= 8'h00;
		14'h0ed6:	ff_dbi <= 8'h00;
		14'h0ed7:	ff_dbi <= 8'h00;
		14'h0ed8:	ff_dbi <= 8'h00;
		14'h0ed9:	ff_dbi <= 8'h00;
		14'h0eda:	ff_dbi <= 8'h00;
		14'h0edb:	ff_dbi <= 8'h00;
		14'h0edc:	ff_dbi <= 8'h00;
		14'h0edd:	ff_dbi <= 8'h00;
		14'h0ede:	ff_dbi <= 8'h00;
		14'h0edf:	ff_dbi <= 8'h00;
		14'h0ee0:	ff_dbi <= 8'h00;
		14'h0ee1:	ff_dbi <= 8'h00;
		14'h0ee2:	ff_dbi <= 8'h00;
		14'h0ee3:	ff_dbi <= 8'h00;
		14'h0ee4:	ff_dbi <= 8'h00;
		14'h0ee5:	ff_dbi <= 8'h00;
		14'h0ee6:	ff_dbi <= 8'h00;
		14'h0ee7:	ff_dbi <= 8'h00;
		14'h0ee8:	ff_dbi <= 8'h00;
		14'h0ee9:	ff_dbi <= 8'h00;
		14'h0eea:	ff_dbi <= 8'h00;
		14'h0eeb:	ff_dbi <= 8'h00;
		14'h0eec:	ff_dbi <= 8'h00;
		14'h0eed:	ff_dbi <= 8'h00;
		14'h0eee:	ff_dbi <= 8'h00;
		14'h0eef:	ff_dbi <= 8'h00;
		14'h0ef0:	ff_dbi <= 8'h00;
		14'h0ef1:	ff_dbi <= 8'h00;
		14'h0ef2:	ff_dbi <= 8'h00;
		14'h0ef3:	ff_dbi <= 8'h00;
		14'h0ef4:	ff_dbi <= 8'h00;
		14'h0ef5:	ff_dbi <= 8'h00;
		14'h0ef6:	ff_dbi <= 8'h00;
		14'h0ef7:	ff_dbi <= 8'h00;
		14'h0ef8:	ff_dbi <= 8'h00;
		14'h0ef9:	ff_dbi <= 8'h00;
		14'h0efa:	ff_dbi <= 8'h00;
		14'h0efb:	ff_dbi <= 8'h00;
		14'h0efc:	ff_dbi <= 8'h00;
		14'h0efd:	ff_dbi <= 8'h00;
		14'h0efe:	ff_dbi <= 8'h00;
		14'h0eff:	ff_dbi <= 8'h00;
		14'h0f00:	ff_dbi <= 8'h00;
		14'h0f01:	ff_dbi <= 8'h00;
		14'h0f02:	ff_dbi <= 8'h00;
		14'h0f03:	ff_dbi <= 8'h00;
		14'h0f04:	ff_dbi <= 8'h00;
		14'h0f05:	ff_dbi <= 8'h00;
		14'h0f06:	ff_dbi <= 8'h00;
		14'h0f07:	ff_dbi <= 8'h00;
		14'h0f08:	ff_dbi <= 8'h00;
		14'h0f09:	ff_dbi <= 8'h00;
		14'h0f0a:	ff_dbi <= 8'h00;
		14'h0f0b:	ff_dbi <= 8'h00;
		14'h0f0c:	ff_dbi <= 8'h00;
		14'h0f0d:	ff_dbi <= 8'h00;
		14'h0f0e:	ff_dbi <= 8'h00;
		14'h0f0f:	ff_dbi <= 8'h00;
		14'h0f10:	ff_dbi <= 8'h00;
		14'h0f11:	ff_dbi <= 8'h00;
		14'h0f12:	ff_dbi <= 8'h00;
		14'h0f13:	ff_dbi <= 8'h00;
		14'h0f14:	ff_dbi <= 8'h00;
		14'h0f15:	ff_dbi <= 8'h00;
		14'h0f16:	ff_dbi <= 8'h00;
		14'h0f17:	ff_dbi <= 8'h00;
		14'h0f18:	ff_dbi <= 8'h00;
		14'h0f19:	ff_dbi <= 8'h00;
		14'h0f1a:	ff_dbi <= 8'h00;
		14'h0f1b:	ff_dbi <= 8'h00;
		14'h0f1c:	ff_dbi <= 8'h00;
		14'h0f1d:	ff_dbi <= 8'h00;
		14'h0f1e:	ff_dbi <= 8'h00;
		14'h0f1f:	ff_dbi <= 8'h00;
		14'h0f20:	ff_dbi <= 8'h00;
		14'h0f21:	ff_dbi <= 8'h00;
		14'h0f22:	ff_dbi <= 8'h00;
		14'h0f23:	ff_dbi <= 8'h00;
		14'h0f24:	ff_dbi <= 8'h00;
		14'h0f25:	ff_dbi <= 8'h00;
		14'h0f26:	ff_dbi <= 8'h00;
		14'h0f27:	ff_dbi <= 8'h00;
		14'h0f28:	ff_dbi <= 8'h00;
		14'h0f29:	ff_dbi <= 8'h00;
		14'h0f2a:	ff_dbi <= 8'h00;
		14'h0f2b:	ff_dbi <= 8'h00;
		14'h0f2c:	ff_dbi <= 8'h00;
		14'h0f2d:	ff_dbi <= 8'h00;
		14'h0f2e:	ff_dbi <= 8'h00;
		14'h0f2f:	ff_dbi <= 8'h00;
		14'h0f30:	ff_dbi <= 8'h00;
		14'h0f31:	ff_dbi <= 8'h00;
		14'h0f32:	ff_dbi <= 8'h00;
		14'h0f33:	ff_dbi <= 8'h00;
		14'h0f34:	ff_dbi <= 8'h00;
		14'h0f35:	ff_dbi <= 8'h00;
		14'h0f36:	ff_dbi <= 8'h00;
		14'h0f37:	ff_dbi <= 8'h00;
		14'h0f38:	ff_dbi <= 8'h00;
		14'h0f39:	ff_dbi <= 8'h00;
		14'h0f3a:	ff_dbi <= 8'h00;
		14'h0f3b:	ff_dbi <= 8'h00;
		14'h0f3c:	ff_dbi <= 8'h00;
		14'h0f3d:	ff_dbi <= 8'h00;
		14'h0f3e:	ff_dbi <= 8'h00;
		14'h0f3f:	ff_dbi <= 8'h00;
		14'h0f40:	ff_dbi <= 8'h00;
		14'h0f41:	ff_dbi <= 8'h00;
		14'h0f42:	ff_dbi <= 8'h00;
		14'h0f43:	ff_dbi <= 8'h00;
		14'h0f44:	ff_dbi <= 8'h00;
		14'h0f45:	ff_dbi <= 8'h00;
		14'h0f46:	ff_dbi <= 8'h00;
		14'h0f47:	ff_dbi <= 8'h00;
		14'h0f48:	ff_dbi <= 8'h00;
		14'h0f49:	ff_dbi <= 8'h00;
		14'h0f4a:	ff_dbi <= 8'h00;
		14'h0f4b:	ff_dbi <= 8'h00;
		14'h0f4c:	ff_dbi <= 8'h00;
		14'h0f4d:	ff_dbi <= 8'h00;
		14'h0f4e:	ff_dbi <= 8'h00;
		14'h0f4f:	ff_dbi <= 8'h00;
		14'h0f50:	ff_dbi <= 8'h00;
		14'h0f51:	ff_dbi <= 8'h00;
		14'h0f52:	ff_dbi <= 8'h00;
		14'h0f53:	ff_dbi <= 8'h00;
		14'h0f54:	ff_dbi <= 8'h00;
		14'h0f55:	ff_dbi <= 8'h00;
		14'h0f56:	ff_dbi <= 8'h00;
		14'h0f57:	ff_dbi <= 8'h00;
		14'h0f58:	ff_dbi <= 8'h00;
		14'h0f59:	ff_dbi <= 8'h00;
		14'h0f5a:	ff_dbi <= 8'h00;
		14'h0f5b:	ff_dbi <= 8'h00;
		14'h0f5c:	ff_dbi <= 8'h00;
		14'h0f5d:	ff_dbi <= 8'h00;
		14'h0f5e:	ff_dbi <= 8'h00;
		14'h0f5f:	ff_dbi <= 8'h00;
		14'h0f60:	ff_dbi <= 8'h00;
		14'h0f61:	ff_dbi <= 8'h00;
		14'h0f62:	ff_dbi <= 8'h00;
		14'h0f63:	ff_dbi <= 8'h00;
		14'h0f64:	ff_dbi <= 8'h00;
		14'h0f65:	ff_dbi <= 8'h00;
		14'h0f66:	ff_dbi <= 8'h00;
		14'h0f67:	ff_dbi <= 8'h00;
		14'h0f68:	ff_dbi <= 8'h00;
		14'h0f69:	ff_dbi <= 8'h00;
		14'h0f6a:	ff_dbi <= 8'h00;
		14'h0f6b:	ff_dbi <= 8'h00;
		14'h0f6c:	ff_dbi <= 8'h00;
		14'h0f6d:	ff_dbi <= 8'h00;
		14'h0f6e:	ff_dbi <= 8'h00;
		14'h0f6f:	ff_dbi <= 8'h00;
		14'h0f70:	ff_dbi <= 8'h00;
		14'h0f71:	ff_dbi <= 8'h00;
		14'h0f72:	ff_dbi <= 8'h00;
		14'h0f73:	ff_dbi <= 8'h00;
		14'h0f74:	ff_dbi <= 8'h00;
		14'h0f75:	ff_dbi <= 8'h00;
		14'h0f76:	ff_dbi <= 8'h00;
		14'h0f77:	ff_dbi <= 8'h00;
		14'h0f78:	ff_dbi <= 8'h00;
		14'h0f79:	ff_dbi <= 8'h00;
		14'h0f7a:	ff_dbi <= 8'h00;
		14'h0f7b:	ff_dbi <= 8'h00;
		14'h0f7c:	ff_dbi <= 8'h00;
		14'h0f7d:	ff_dbi <= 8'h00;
		14'h0f7e:	ff_dbi <= 8'h00;
		14'h0f7f:	ff_dbi <= 8'h00;
		14'h0f80:	ff_dbi <= 8'h00;
		14'h0f81:	ff_dbi <= 8'h00;
		14'h0f82:	ff_dbi <= 8'h00;
		14'h0f83:	ff_dbi <= 8'h00;
		14'h0f84:	ff_dbi <= 8'h00;
		14'h0f85:	ff_dbi <= 8'h00;
		14'h0f86:	ff_dbi <= 8'h00;
		14'h0f87:	ff_dbi <= 8'h00;
		14'h0f88:	ff_dbi <= 8'h00;
		14'h0f89:	ff_dbi <= 8'h00;
		14'h0f8a:	ff_dbi <= 8'h00;
		14'h0f8b:	ff_dbi <= 8'h00;
		14'h0f8c:	ff_dbi <= 8'h00;
		14'h0f8d:	ff_dbi <= 8'h00;
		14'h0f8e:	ff_dbi <= 8'h00;
		14'h0f8f:	ff_dbi <= 8'h00;
		14'h0f90:	ff_dbi <= 8'h00;
		14'h0f91:	ff_dbi <= 8'h00;
		14'h0f92:	ff_dbi <= 8'h00;
		14'h0f93:	ff_dbi <= 8'h00;
		14'h0f94:	ff_dbi <= 8'h00;
		14'h0f95:	ff_dbi <= 8'h00;
		14'h0f96:	ff_dbi <= 8'h00;
		14'h0f97:	ff_dbi <= 8'h00;
		14'h0f98:	ff_dbi <= 8'h00;
		14'h0f99:	ff_dbi <= 8'h00;
		14'h0f9a:	ff_dbi <= 8'h00;
		14'h0f9b:	ff_dbi <= 8'h00;
		14'h0f9c:	ff_dbi <= 8'h00;
		14'h0f9d:	ff_dbi <= 8'h00;
		14'h0f9e:	ff_dbi <= 8'h00;
		14'h0f9f:	ff_dbi <= 8'h00;
		14'h0fa0:	ff_dbi <= 8'h00;
		14'h0fa1:	ff_dbi <= 8'h00;
		14'h0fa2:	ff_dbi <= 8'h00;
		14'h0fa3:	ff_dbi <= 8'h00;
		14'h0fa4:	ff_dbi <= 8'h00;
		14'h0fa5:	ff_dbi <= 8'h00;
		14'h0fa6:	ff_dbi <= 8'h00;
		14'h0fa7:	ff_dbi <= 8'h00;
		14'h0fa8:	ff_dbi <= 8'h00;
		14'h0fa9:	ff_dbi <= 8'h00;
		14'h0faa:	ff_dbi <= 8'h00;
		14'h0fab:	ff_dbi <= 8'h00;
		14'h0fac:	ff_dbi <= 8'h00;
		14'h0fad:	ff_dbi <= 8'h00;
		14'h0fae:	ff_dbi <= 8'h00;
		14'h0faf:	ff_dbi <= 8'h00;
		14'h0fb0:	ff_dbi <= 8'h00;
		14'h0fb1:	ff_dbi <= 8'h00;
		14'h0fb2:	ff_dbi <= 8'h00;
		14'h0fb3:	ff_dbi <= 8'h00;
		14'h0fb4:	ff_dbi <= 8'h00;
		14'h0fb5:	ff_dbi <= 8'h00;
		14'h0fb6:	ff_dbi <= 8'h00;
		14'h0fb7:	ff_dbi <= 8'h00;
		14'h0fb8:	ff_dbi <= 8'h00;
		14'h0fb9:	ff_dbi <= 8'h00;
		14'h0fba:	ff_dbi <= 8'h00;
		14'h0fbb:	ff_dbi <= 8'h00;
		14'h0fbc:	ff_dbi <= 8'h00;
		14'h0fbd:	ff_dbi <= 8'h00;
		14'h0fbe:	ff_dbi <= 8'h00;
		14'h0fbf:	ff_dbi <= 8'h00;
		14'h0fc0:	ff_dbi <= 8'h00;
		14'h0fc1:	ff_dbi <= 8'h00;
		14'h0fc2:	ff_dbi <= 8'h00;
		14'h0fc3:	ff_dbi <= 8'h00;
		14'h0fc4:	ff_dbi <= 8'h00;
		14'h0fc5:	ff_dbi <= 8'h00;
		14'h0fc6:	ff_dbi <= 8'h00;
		14'h0fc7:	ff_dbi <= 8'h00;
		14'h0fc8:	ff_dbi <= 8'h00;
		14'h0fc9:	ff_dbi <= 8'h00;
		14'h0fca:	ff_dbi <= 8'h00;
		14'h0fcb:	ff_dbi <= 8'h00;
		14'h0fcc:	ff_dbi <= 8'h00;
		14'h0fcd:	ff_dbi <= 8'h00;
		14'h0fce:	ff_dbi <= 8'h00;
		14'h0fcf:	ff_dbi <= 8'h00;
		14'h0fd0:	ff_dbi <= 8'h00;
		14'h0fd1:	ff_dbi <= 8'h00;
		14'h0fd2:	ff_dbi <= 8'h00;
		14'h0fd3:	ff_dbi <= 8'h00;
		14'h0fd4:	ff_dbi <= 8'h00;
		14'h0fd5:	ff_dbi <= 8'h00;
		14'h0fd6:	ff_dbi <= 8'h00;
		14'h0fd7:	ff_dbi <= 8'h00;
		14'h0fd8:	ff_dbi <= 8'h00;
		14'h0fd9:	ff_dbi <= 8'h00;
		14'h0fda:	ff_dbi <= 8'h00;
		14'h0fdb:	ff_dbi <= 8'h00;
		14'h0fdc:	ff_dbi <= 8'h00;
		14'h0fdd:	ff_dbi <= 8'h00;
		14'h0fde:	ff_dbi <= 8'h00;
		14'h0fdf:	ff_dbi <= 8'h00;
		14'h0fe0:	ff_dbi <= 8'h00;
		14'h0fe1:	ff_dbi <= 8'h00;
		14'h0fe2:	ff_dbi <= 8'h00;
		14'h0fe3:	ff_dbi <= 8'h00;
		14'h0fe4:	ff_dbi <= 8'h00;
		14'h0fe5:	ff_dbi <= 8'h00;
		14'h0fe6:	ff_dbi <= 8'h00;
		14'h0fe7:	ff_dbi <= 8'h00;
		14'h0fe8:	ff_dbi <= 8'h00;
		14'h0fe9:	ff_dbi <= 8'h00;
		14'h0fea:	ff_dbi <= 8'h00;
		14'h0feb:	ff_dbi <= 8'h00;
		14'h0fec:	ff_dbi <= 8'h00;
		14'h0fed:	ff_dbi <= 8'h00;
		14'h0fee:	ff_dbi <= 8'h00;
		14'h0fef:	ff_dbi <= 8'h00;
		14'h0ff0:	ff_dbi <= 8'h00;
		14'h0ff1:	ff_dbi <= 8'h00;
		14'h0ff2:	ff_dbi <= 8'h00;
		14'h0ff3:	ff_dbi <= 8'h00;
		14'h0ff4:	ff_dbi <= 8'h00;
		14'h0ff5:	ff_dbi <= 8'h00;
		14'h0ff6:	ff_dbi <= 8'h00;
		14'h0ff7:	ff_dbi <= 8'h00;
		14'h0ff8:	ff_dbi <= 8'h00;
		14'h0ff9:	ff_dbi <= 8'h00;
		14'h0ffa:	ff_dbi <= 8'h00;
		14'h0ffb:	ff_dbi <= 8'h00;
		14'h0ffc:	ff_dbi <= 8'h00;
		14'h0ffd:	ff_dbi <= 8'h00;
		14'h0ffe:	ff_dbi <= 8'h00;
		14'h0fff:	ff_dbi <= 8'h00;
		14'h1000:	ff_dbi <= 8'h00;
		14'h1001:	ff_dbi <= 8'h00;
		14'h1002:	ff_dbi <= 8'h00;
		14'h1003:	ff_dbi <= 8'h00;
		14'h1004:	ff_dbi <= 8'h00;
		14'h1005:	ff_dbi <= 8'h00;
		14'h1006:	ff_dbi <= 8'h00;
		14'h1007:	ff_dbi <= 8'h00;
		14'h1008:	ff_dbi <= 8'h00;
		14'h1009:	ff_dbi <= 8'h00;
		14'h100a:	ff_dbi <= 8'h00;
		14'h100b:	ff_dbi <= 8'h00;
		14'h100c:	ff_dbi <= 8'h00;
		14'h100d:	ff_dbi <= 8'h00;
		14'h100e:	ff_dbi <= 8'h00;
		14'h100f:	ff_dbi <= 8'h00;
		14'h1010:	ff_dbi <= 8'h00;
		14'h1011:	ff_dbi <= 8'h00;
		14'h1012:	ff_dbi <= 8'h00;
		14'h1013:	ff_dbi <= 8'h00;
		14'h1014:	ff_dbi <= 8'h00;
		14'h1015:	ff_dbi <= 8'h00;
		14'h1016:	ff_dbi <= 8'h00;
		14'h1017:	ff_dbi <= 8'h00;
		14'h1018:	ff_dbi <= 8'h00;
		14'h1019:	ff_dbi <= 8'h00;
		14'h101a:	ff_dbi <= 8'h00;
		14'h101b:	ff_dbi <= 8'h00;
		14'h101c:	ff_dbi <= 8'h00;
		14'h101d:	ff_dbi <= 8'h00;
		14'h101e:	ff_dbi <= 8'h00;
		14'h101f:	ff_dbi <= 8'h00;
		14'h1020:	ff_dbi <= 8'h00;
		14'h1021:	ff_dbi <= 8'h00;
		14'h1022:	ff_dbi <= 8'h00;
		14'h1023:	ff_dbi <= 8'h00;
		14'h1024:	ff_dbi <= 8'h00;
		14'h1025:	ff_dbi <= 8'h00;
		14'h1026:	ff_dbi <= 8'h00;
		14'h1027:	ff_dbi <= 8'h00;
		14'h1028:	ff_dbi <= 8'h00;
		14'h1029:	ff_dbi <= 8'h00;
		14'h102a:	ff_dbi <= 8'h00;
		14'h102b:	ff_dbi <= 8'h00;
		14'h102c:	ff_dbi <= 8'h00;
		14'h102d:	ff_dbi <= 8'h00;
		14'h102e:	ff_dbi <= 8'h00;
		14'h102f:	ff_dbi <= 8'h00;
		14'h1030:	ff_dbi <= 8'h00;
		14'h1031:	ff_dbi <= 8'h00;
		14'h1032:	ff_dbi <= 8'h00;
		14'h1033:	ff_dbi <= 8'h00;
		14'h1034:	ff_dbi <= 8'h00;
		14'h1035:	ff_dbi <= 8'h00;
		14'h1036:	ff_dbi <= 8'h00;
		14'h1037:	ff_dbi <= 8'h00;
		14'h1038:	ff_dbi <= 8'h00;
		14'h1039:	ff_dbi <= 8'h00;
		14'h103a:	ff_dbi <= 8'h00;
		14'h103b:	ff_dbi <= 8'h00;
		14'h103c:	ff_dbi <= 8'h00;
		14'h103d:	ff_dbi <= 8'h00;
		14'h103e:	ff_dbi <= 8'h00;
		14'h103f:	ff_dbi <= 8'h00;
		14'h1040:	ff_dbi <= 8'h00;
		14'h1041:	ff_dbi <= 8'h00;
		14'h1042:	ff_dbi <= 8'h00;
		14'h1043:	ff_dbi <= 8'h00;
		14'h1044:	ff_dbi <= 8'h00;
		14'h1045:	ff_dbi <= 8'h00;
		14'h1046:	ff_dbi <= 8'h00;
		14'h1047:	ff_dbi <= 8'h00;
		14'h1048:	ff_dbi <= 8'h00;
		14'h1049:	ff_dbi <= 8'h00;
		14'h104a:	ff_dbi <= 8'h00;
		14'h104b:	ff_dbi <= 8'h00;
		14'h104c:	ff_dbi <= 8'h00;
		14'h104d:	ff_dbi <= 8'h00;
		14'h104e:	ff_dbi <= 8'h00;
		14'h104f:	ff_dbi <= 8'h00;
		14'h1050:	ff_dbi <= 8'h00;
		14'h1051:	ff_dbi <= 8'h00;
		14'h1052:	ff_dbi <= 8'h00;
		14'h1053:	ff_dbi <= 8'h00;
		14'h1054:	ff_dbi <= 8'h00;
		14'h1055:	ff_dbi <= 8'h00;
		14'h1056:	ff_dbi <= 8'h00;
		14'h1057:	ff_dbi <= 8'h00;
		14'h1058:	ff_dbi <= 8'h00;
		14'h1059:	ff_dbi <= 8'h00;
		14'h105a:	ff_dbi <= 8'h00;
		14'h105b:	ff_dbi <= 8'h00;
		14'h105c:	ff_dbi <= 8'h00;
		14'h105d:	ff_dbi <= 8'h00;
		14'h105e:	ff_dbi <= 8'h00;
		14'h105f:	ff_dbi <= 8'h00;
		14'h1060:	ff_dbi <= 8'h00;
		14'h1061:	ff_dbi <= 8'h00;
		14'h1062:	ff_dbi <= 8'h00;
		14'h1063:	ff_dbi <= 8'h00;
		14'h1064:	ff_dbi <= 8'h00;
		14'h1065:	ff_dbi <= 8'h00;
		14'h1066:	ff_dbi <= 8'h00;
		14'h1067:	ff_dbi <= 8'h00;
		14'h1068:	ff_dbi <= 8'h00;
		14'h1069:	ff_dbi <= 8'h00;
		14'h106a:	ff_dbi <= 8'h00;
		14'h106b:	ff_dbi <= 8'h00;
		14'h106c:	ff_dbi <= 8'h00;
		14'h106d:	ff_dbi <= 8'h00;
		14'h106e:	ff_dbi <= 8'h00;
		14'h106f:	ff_dbi <= 8'h00;
		14'h1070:	ff_dbi <= 8'h00;
		14'h1071:	ff_dbi <= 8'h00;
		14'h1072:	ff_dbi <= 8'h00;
		14'h1073:	ff_dbi <= 8'h00;
		14'h1074:	ff_dbi <= 8'h00;
		14'h1075:	ff_dbi <= 8'h00;
		14'h1076:	ff_dbi <= 8'h00;
		14'h1077:	ff_dbi <= 8'h00;
		14'h1078:	ff_dbi <= 8'h00;
		14'h1079:	ff_dbi <= 8'h00;
		14'h107a:	ff_dbi <= 8'h00;
		14'h107b:	ff_dbi <= 8'h00;
		14'h107c:	ff_dbi <= 8'h00;
		14'h107d:	ff_dbi <= 8'h00;
		14'h107e:	ff_dbi <= 8'h00;
		14'h107f:	ff_dbi <= 8'h00;
		14'h1080:	ff_dbi <= 8'h00;
		14'h1081:	ff_dbi <= 8'h00;
		14'h1082:	ff_dbi <= 8'h00;
		14'h1083:	ff_dbi <= 8'h00;
		14'h1084:	ff_dbi <= 8'h00;
		14'h1085:	ff_dbi <= 8'h00;
		14'h1086:	ff_dbi <= 8'h00;
		14'h1087:	ff_dbi <= 8'h00;
		14'h1088:	ff_dbi <= 8'h00;
		14'h1089:	ff_dbi <= 8'h00;
		14'h108a:	ff_dbi <= 8'h00;
		14'h108b:	ff_dbi <= 8'h00;
		14'h108c:	ff_dbi <= 8'h00;
		14'h108d:	ff_dbi <= 8'h00;
		14'h108e:	ff_dbi <= 8'h00;
		14'h108f:	ff_dbi <= 8'h00;
		14'h1090:	ff_dbi <= 8'h00;
		14'h1091:	ff_dbi <= 8'h00;
		14'h1092:	ff_dbi <= 8'h00;
		14'h1093:	ff_dbi <= 8'h00;
		14'h1094:	ff_dbi <= 8'h00;
		14'h1095:	ff_dbi <= 8'h00;
		14'h1096:	ff_dbi <= 8'h00;
		14'h1097:	ff_dbi <= 8'h00;
		14'h1098:	ff_dbi <= 8'h00;
		14'h1099:	ff_dbi <= 8'h00;
		14'h109a:	ff_dbi <= 8'h00;
		14'h109b:	ff_dbi <= 8'h00;
		14'h109c:	ff_dbi <= 8'h00;
		14'h109d:	ff_dbi <= 8'h00;
		14'h109e:	ff_dbi <= 8'h00;
		14'h109f:	ff_dbi <= 8'h00;
		14'h10a0:	ff_dbi <= 8'h00;
		14'h10a1:	ff_dbi <= 8'h00;
		14'h10a2:	ff_dbi <= 8'h00;
		14'h10a3:	ff_dbi <= 8'h00;
		14'h10a4:	ff_dbi <= 8'h00;
		14'h10a5:	ff_dbi <= 8'h00;
		14'h10a6:	ff_dbi <= 8'h00;
		14'h10a7:	ff_dbi <= 8'h00;
		14'h10a8:	ff_dbi <= 8'h00;
		14'h10a9:	ff_dbi <= 8'h00;
		14'h10aa:	ff_dbi <= 8'h00;
		14'h10ab:	ff_dbi <= 8'h00;
		14'h10ac:	ff_dbi <= 8'h00;
		14'h10ad:	ff_dbi <= 8'h00;
		14'h10ae:	ff_dbi <= 8'h00;
		14'h10af:	ff_dbi <= 8'h00;
		14'h10b0:	ff_dbi <= 8'h00;
		14'h10b1:	ff_dbi <= 8'h00;
		14'h10b2:	ff_dbi <= 8'h00;
		14'h10b3:	ff_dbi <= 8'h00;
		14'h10b4:	ff_dbi <= 8'h00;
		14'h10b5:	ff_dbi <= 8'h00;
		14'h10b6:	ff_dbi <= 8'h00;
		14'h10b7:	ff_dbi <= 8'h00;
		14'h10b8:	ff_dbi <= 8'h00;
		14'h10b9:	ff_dbi <= 8'h00;
		14'h10ba:	ff_dbi <= 8'h00;
		14'h10bb:	ff_dbi <= 8'h00;
		14'h10bc:	ff_dbi <= 8'h00;
		14'h10bd:	ff_dbi <= 8'h00;
		14'h10be:	ff_dbi <= 8'h00;
		14'h10bf:	ff_dbi <= 8'h00;
		14'h10c0:	ff_dbi <= 8'h00;
		14'h10c1:	ff_dbi <= 8'h00;
		14'h10c2:	ff_dbi <= 8'h00;
		14'h10c3:	ff_dbi <= 8'h00;
		14'h10c4:	ff_dbi <= 8'h00;
		14'h10c5:	ff_dbi <= 8'h00;
		14'h10c6:	ff_dbi <= 8'h00;
		14'h10c7:	ff_dbi <= 8'h00;
		14'h10c8:	ff_dbi <= 8'h00;
		14'h10c9:	ff_dbi <= 8'h00;
		14'h10ca:	ff_dbi <= 8'h00;
		14'h10cb:	ff_dbi <= 8'h00;
		14'h10cc:	ff_dbi <= 8'h00;
		14'h10cd:	ff_dbi <= 8'h00;
		14'h10ce:	ff_dbi <= 8'h00;
		14'h10cf:	ff_dbi <= 8'h00;
		14'h10d0:	ff_dbi <= 8'h00;
		14'h10d1:	ff_dbi <= 8'h00;
		14'h10d2:	ff_dbi <= 8'h00;
		14'h10d3:	ff_dbi <= 8'h00;
		14'h10d4:	ff_dbi <= 8'h00;
		14'h10d5:	ff_dbi <= 8'h00;
		14'h10d6:	ff_dbi <= 8'h00;
		14'h10d7:	ff_dbi <= 8'h00;
		14'h10d8:	ff_dbi <= 8'h00;
		14'h10d9:	ff_dbi <= 8'h00;
		14'h10da:	ff_dbi <= 8'h00;
		14'h10db:	ff_dbi <= 8'h00;
		14'h10dc:	ff_dbi <= 8'h00;
		14'h10dd:	ff_dbi <= 8'h00;
		14'h10de:	ff_dbi <= 8'h00;
		14'h10df:	ff_dbi <= 8'h00;
		14'h10e0:	ff_dbi <= 8'h00;
		14'h10e1:	ff_dbi <= 8'h00;
		14'h10e2:	ff_dbi <= 8'h00;
		14'h10e3:	ff_dbi <= 8'h00;
		14'h10e4:	ff_dbi <= 8'h00;
		14'h10e5:	ff_dbi <= 8'h00;
		14'h10e6:	ff_dbi <= 8'h00;
		14'h10e7:	ff_dbi <= 8'h00;
		14'h10e8:	ff_dbi <= 8'h00;
		14'h10e9:	ff_dbi <= 8'h00;
		14'h10ea:	ff_dbi <= 8'h00;
		14'h10eb:	ff_dbi <= 8'h00;
		14'h10ec:	ff_dbi <= 8'h00;
		14'h10ed:	ff_dbi <= 8'h00;
		14'h10ee:	ff_dbi <= 8'h00;
		14'h10ef:	ff_dbi <= 8'h00;
		14'h10f0:	ff_dbi <= 8'h00;
		14'h10f1:	ff_dbi <= 8'h00;
		14'h10f2:	ff_dbi <= 8'h00;
		14'h10f3:	ff_dbi <= 8'h00;
		14'h10f4:	ff_dbi <= 8'h00;
		14'h10f5:	ff_dbi <= 8'h00;
		14'h10f6:	ff_dbi <= 8'h00;
		14'h10f7:	ff_dbi <= 8'h00;
		14'h10f8:	ff_dbi <= 8'h00;
		14'h10f9:	ff_dbi <= 8'h00;
		14'h10fa:	ff_dbi <= 8'h00;
		14'h10fb:	ff_dbi <= 8'h00;
		14'h10fc:	ff_dbi <= 8'h00;
		14'h10fd:	ff_dbi <= 8'h00;
		14'h10fe:	ff_dbi <= 8'h00;
		14'h10ff:	ff_dbi <= 8'h00;
		14'h1100:	ff_dbi <= 8'h00;
		14'h1101:	ff_dbi <= 8'h00;
		14'h1102:	ff_dbi <= 8'h00;
		14'h1103:	ff_dbi <= 8'h00;
		14'h1104:	ff_dbi <= 8'h00;
		14'h1105:	ff_dbi <= 8'h00;
		14'h1106:	ff_dbi <= 8'h00;
		14'h1107:	ff_dbi <= 8'h00;
		14'h1108:	ff_dbi <= 8'h00;
		14'h1109:	ff_dbi <= 8'h00;
		14'h110a:	ff_dbi <= 8'h00;
		14'h110b:	ff_dbi <= 8'h00;
		14'h110c:	ff_dbi <= 8'h00;
		14'h110d:	ff_dbi <= 8'h00;
		14'h110e:	ff_dbi <= 8'h00;
		14'h110f:	ff_dbi <= 8'h00;
		14'h1110:	ff_dbi <= 8'h00;
		14'h1111:	ff_dbi <= 8'h00;
		14'h1112:	ff_dbi <= 8'h00;
		14'h1113:	ff_dbi <= 8'h00;
		14'h1114:	ff_dbi <= 8'h00;
		14'h1115:	ff_dbi <= 8'h00;
		14'h1116:	ff_dbi <= 8'h00;
		14'h1117:	ff_dbi <= 8'h00;
		14'h1118:	ff_dbi <= 8'h00;
		14'h1119:	ff_dbi <= 8'h00;
		14'h111a:	ff_dbi <= 8'h00;
		14'h111b:	ff_dbi <= 8'h00;
		14'h111c:	ff_dbi <= 8'h00;
		14'h111d:	ff_dbi <= 8'h00;
		14'h111e:	ff_dbi <= 8'h00;
		14'h111f:	ff_dbi <= 8'h00;
		14'h1120:	ff_dbi <= 8'h00;
		14'h1121:	ff_dbi <= 8'h00;
		14'h1122:	ff_dbi <= 8'h00;
		14'h1123:	ff_dbi <= 8'h00;
		14'h1124:	ff_dbi <= 8'h00;
		14'h1125:	ff_dbi <= 8'h00;
		14'h1126:	ff_dbi <= 8'h00;
		14'h1127:	ff_dbi <= 8'h00;
		14'h1128:	ff_dbi <= 8'h00;
		14'h1129:	ff_dbi <= 8'h00;
		14'h112a:	ff_dbi <= 8'h00;
		14'h112b:	ff_dbi <= 8'h00;
		14'h112c:	ff_dbi <= 8'h00;
		14'h112d:	ff_dbi <= 8'h00;
		14'h112e:	ff_dbi <= 8'h00;
		14'h112f:	ff_dbi <= 8'h00;
		14'h1130:	ff_dbi <= 8'h00;
		14'h1131:	ff_dbi <= 8'h00;
		14'h1132:	ff_dbi <= 8'h00;
		14'h1133:	ff_dbi <= 8'h00;
		14'h1134:	ff_dbi <= 8'h00;
		14'h1135:	ff_dbi <= 8'h00;
		14'h1136:	ff_dbi <= 8'h00;
		14'h1137:	ff_dbi <= 8'h00;
		14'h1138:	ff_dbi <= 8'h00;
		14'h1139:	ff_dbi <= 8'h00;
		14'h113a:	ff_dbi <= 8'h00;
		14'h113b:	ff_dbi <= 8'h00;
		14'h113c:	ff_dbi <= 8'h00;
		14'h113d:	ff_dbi <= 8'h00;
		14'h113e:	ff_dbi <= 8'h00;
		14'h113f:	ff_dbi <= 8'h00;
		14'h1140:	ff_dbi <= 8'h00;
		14'h1141:	ff_dbi <= 8'h00;
		14'h1142:	ff_dbi <= 8'h00;
		14'h1143:	ff_dbi <= 8'h00;
		14'h1144:	ff_dbi <= 8'h00;
		14'h1145:	ff_dbi <= 8'h00;
		14'h1146:	ff_dbi <= 8'h00;
		14'h1147:	ff_dbi <= 8'h00;
		14'h1148:	ff_dbi <= 8'h00;
		14'h1149:	ff_dbi <= 8'h00;
		14'h114a:	ff_dbi <= 8'h00;
		14'h114b:	ff_dbi <= 8'h00;
		14'h114c:	ff_dbi <= 8'h00;
		14'h114d:	ff_dbi <= 8'h00;
		14'h114e:	ff_dbi <= 8'h00;
		14'h114f:	ff_dbi <= 8'h00;
		14'h1150:	ff_dbi <= 8'h00;
		14'h1151:	ff_dbi <= 8'h00;
		14'h1152:	ff_dbi <= 8'h00;
		14'h1153:	ff_dbi <= 8'h00;
		14'h1154:	ff_dbi <= 8'h00;
		14'h1155:	ff_dbi <= 8'h00;
		14'h1156:	ff_dbi <= 8'h00;
		14'h1157:	ff_dbi <= 8'h00;
		14'h1158:	ff_dbi <= 8'h00;
		14'h1159:	ff_dbi <= 8'h00;
		14'h115a:	ff_dbi <= 8'h00;
		14'h115b:	ff_dbi <= 8'h00;
		14'h115c:	ff_dbi <= 8'h00;
		14'h115d:	ff_dbi <= 8'h00;
		14'h115e:	ff_dbi <= 8'h00;
		14'h115f:	ff_dbi <= 8'h00;
		14'h1160:	ff_dbi <= 8'h00;
		14'h1161:	ff_dbi <= 8'h00;
		14'h1162:	ff_dbi <= 8'h00;
		14'h1163:	ff_dbi <= 8'h00;
		14'h1164:	ff_dbi <= 8'h00;
		14'h1165:	ff_dbi <= 8'h00;
		14'h1166:	ff_dbi <= 8'h00;
		14'h1167:	ff_dbi <= 8'h00;
		14'h1168:	ff_dbi <= 8'h00;
		14'h1169:	ff_dbi <= 8'h00;
		14'h116a:	ff_dbi <= 8'h00;
		14'h116b:	ff_dbi <= 8'h00;
		14'h116c:	ff_dbi <= 8'h00;
		14'h116d:	ff_dbi <= 8'h00;
		14'h116e:	ff_dbi <= 8'h00;
		14'h116f:	ff_dbi <= 8'h00;
		14'h1170:	ff_dbi <= 8'h00;
		14'h1171:	ff_dbi <= 8'h00;
		14'h1172:	ff_dbi <= 8'h00;
		14'h1173:	ff_dbi <= 8'h00;
		14'h1174:	ff_dbi <= 8'h00;
		14'h1175:	ff_dbi <= 8'h00;
		14'h1176:	ff_dbi <= 8'h00;
		14'h1177:	ff_dbi <= 8'h00;
		14'h1178:	ff_dbi <= 8'h00;
		14'h1179:	ff_dbi <= 8'h00;
		14'h117a:	ff_dbi <= 8'h00;
		14'h117b:	ff_dbi <= 8'h00;
		14'h117c:	ff_dbi <= 8'h00;
		14'h117d:	ff_dbi <= 8'h00;
		14'h117e:	ff_dbi <= 8'h00;
		14'h117f:	ff_dbi <= 8'h00;
		14'h1180:	ff_dbi <= 8'h00;
		14'h1181:	ff_dbi <= 8'h00;
		14'h1182:	ff_dbi <= 8'h00;
		14'h1183:	ff_dbi <= 8'h00;
		14'h1184:	ff_dbi <= 8'h00;
		14'h1185:	ff_dbi <= 8'h00;
		14'h1186:	ff_dbi <= 8'h00;
		14'h1187:	ff_dbi <= 8'h00;
		14'h1188:	ff_dbi <= 8'h00;
		14'h1189:	ff_dbi <= 8'h00;
		14'h118a:	ff_dbi <= 8'h00;
		14'h118b:	ff_dbi <= 8'h00;
		14'h118c:	ff_dbi <= 8'h00;
		14'h118d:	ff_dbi <= 8'h00;
		14'h118e:	ff_dbi <= 8'h00;
		14'h118f:	ff_dbi <= 8'h00;
		14'h1190:	ff_dbi <= 8'h00;
		14'h1191:	ff_dbi <= 8'h00;
		14'h1192:	ff_dbi <= 8'h00;
		14'h1193:	ff_dbi <= 8'h00;
		14'h1194:	ff_dbi <= 8'h00;
		14'h1195:	ff_dbi <= 8'h00;
		14'h1196:	ff_dbi <= 8'h00;
		14'h1197:	ff_dbi <= 8'h00;
		14'h1198:	ff_dbi <= 8'h00;
		14'h1199:	ff_dbi <= 8'h00;
		14'h119a:	ff_dbi <= 8'h00;
		14'h119b:	ff_dbi <= 8'h00;
		14'h119c:	ff_dbi <= 8'h00;
		14'h119d:	ff_dbi <= 8'h00;
		14'h119e:	ff_dbi <= 8'h00;
		14'h119f:	ff_dbi <= 8'h00;
		14'h11a0:	ff_dbi <= 8'h00;
		14'h11a1:	ff_dbi <= 8'h00;
		14'h11a2:	ff_dbi <= 8'h00;
		14'h11a3:	ff_dbi <= 8'h00;
		14'h11a4:	ff_dbi <= 8'h00;
		14'h11a5:	ff_dbi <= 8'h00;
		14'h11a6:	ff_dbi <= 8'h00;
		14'h11a7:	ff_dbi <= 8'h00;
		14'h11a8:	ff_dbi <= 8'h00;
		14'h11a9:	ff_dbi <= 8'h00;
		14'h11aa:	ff_dbi <= 8'h00;
		14'h11ab:	ff_dbi <= 8'h00;
		14'h11ac:	ff_dbi <= 8'h00;
		14'h11ad:	ff_dbi <= 8'h00;
		14'h11ae:	ff_dbi <= 8'h00;
		14'h11af:	ff_dbi <= 8'h00;
		14'h11b0:	ff_dbi <= 8'h00;
		14'h11b1:	ff_dbi <= 8'h00;
		14'h11b2:	ff_dbi <= 8'h00;
		14'h11b3:	ff_dbi <= 8'h00;
		14'h11b4:	ff_dbi <= 8'h00;
		14'h11b5:	ff_dbi <= 8'h00;
		14'h11b6:	ff_dbi <= 8'h00;
		14'h11b7:	ff_dbi <= 8'h00;
		14'h11b8:	ff_dbi <= 8'h00;
		14'h11b9:	ff_dbi <= 8'h00;
		14'h11ba:	ff_dbi <= 8'h00;
		14'h11bb:	ff_dbi <= 8'h00;
		14'h11bc:	ff_dbi <= 8'h00;
		14'h11bd:	ff_dbi <= 8'h00;
		14'h11be:	ff_dbi <= 8'h00;
		14'h11bf:	ff_dbi <= 8'h00;
		14'h11c0:	ff_dbi <= 8'h00;
		14'h11c1:	ff_dbi <= 8'h00;
		14'h11c2:	ff_dbi <= 8'h00;
		14'h11c3:	ff_dbi <= 8'h00;
		14'h11c4:	ff_dbi <= 8'h00;
		14'h11c5:	ff_dbi <= 8'h00;
		14'h11c6:	ff_dbi <= 8'h00;
		14'h11c7:	ff_dbi <= 8'h00;
		14'h11c8:	ff_dbi <= 8'h00;
		14'h11c9:	ff_dbi <= 8'h00;
		14'h11ca:	ff_dbi <= 8'h00;
		14'h11cb:	ff_dbi <= 8'h00;
		14'h11cc:	ff_dbi <= 8'h00;
		14'h11cd:	ff_dbi <= 8'h00;
		14'h11ce:	ff_dbi <= 8'h00;
		14'h11cf:	ff_dbi <= 8'h00;
		14'h11d0:	ff_dbi <= 8'h00;
		14'h11d1:	ff_dbi <= 8'h00;
		14'h11d2:	ff_dbi <= 8'h00;
		14'h11d3:	ff_dbi <= 8'h00;
		14'h11d4:	ff_dbi <= 8'h00;
		14'h11d5:	ff_dbi <= 8'h00;
		14'h11d6:	ff_dbi <= 8'h00;
		14'h11d7:	ff_dbi <= 8'h00;
		14'h11d8:	ff_dbi <= 8'h00;
		14'h11d9:	ff_dbi <= 8'h00;
		14'h11da:	ff_dbi <= 8'h00;
		14'h11db:	ff_dbi <= 8'h00;
		14'h11dc:	ff_dbi <= 8'h00;
		14'h11dd:	ff_dbi <= 8'h00;
		14'h11de:	ff_dbi <= 8'h00;
		14'h11df:	ff_dbi <= 8'h00;
		14'h11e0:	ff_dbi <= 8'h00;
		14'h11e1:	ff_dbi <= 8'h00;
		14'h11e2:	ff_dbi <= 8'h00;
		14'h11e3:	ff_dbi <= 8'h00;
		14'h11e4:	ff_dbi <= 8'h00;
		14'h11e5:	ff_dbi <= 8'h00;
		14'h11e6:	ff_dbi <= 8'h00;
		14'h11e7:	ff_dbi <= 8'h00;
		14'h11e8:	ff_dbi <= 8'h00;
		14'h11e9:	ff_dbi <= 8'h00;
		14'h11ea:	ff_dbi <= 8'h00;
		14'h11eb:	ff_dbi <= 8'h00;
		14'h11ec:	ff_dbi <= 8'h00;
		14'h11ed:	ff_dbi <= 8'h00;
		14'h11ee:	ff_dbi <= 8'h00;
		14'h11ef:	ff_dbi <= 8'h00;
		14'h11f0:	ff_dbi <= 8'h00;
		14'h11f1:	ff_dbi <= 8'h00;
		14'h11f2:	ff_dbi <= 8'h00;
		14'h11f3:	ff_dbi <= 8'h00;
		14'h11f4:	ff_dbi <= 8'h00;
		14'h11f5:	ff_dbi <= 8'h00;
		14'h11f6:	ff_dbi <= 8'h00;
		14'h11f7:	ff_dbi <= 8'h00;
		14'h11f8:	ff_dbi <= 8'h00;
		14'h11f9:	ff_dbi <= 8'h00;
		14'h11fa:	ff_dbi <= 8'h00;
		14'h11fb:	ff_dbi <= 8'h00;
		14'h11fc:	ff_dbi <= 8'h00;
		14'h11fd:	ff_dbi <= 8'h00;
		14'h11fe:	ff_dbi <= 8'h00;
		14'h11ff:	ff_dbi <= 8'h00;
		14'h1200:	ff_dbi <= 8'h00;
		14'h1201:	ff_dbi <= 8'h00;
		14'h1202:	ff_dbi <= 8'h00;
		14'h1203:	ff_dbi <= 8'h00;
		14'h1204:	ff_dbi <= 8'h00;
		14'h1205:	ff_dbi <= 8'h00;
		14'h1206:	ff_dbi <= 8'h00;
		14'h1207:	ff_dbi <= 8'h00;
		14'h1208:	ff_dbi <= 8'h00;
		14'h1209:	ff_dbi <= 8'h00;
		14'h120a:	ff_dbi <= 8'h00;
		14'h120b:	ff_dbi <= 8'h00;
		14'h120c:	ff_dbi <= 8'h00;
		14'h120d:	ff_dbi <= 8'h00;
		14'h120e:	ff_dbi <= 8'h00;
		14'h120f:	ff_dbi <= 8'h00;
		14'h1210:	ff_dbi <= 8'h00;
		14'h1211:	ff_dbi <= 8'h00;
		14'h1212:	ff_dbi <= 8'h00;
		14'h1213:	ff_dbi <= 8'h00;
		14'h1214:	ff_dbi <= 8'h00;
		14'h1215:	ff_dbi <= 8'h00;
		14'h1216:	ff_dbi <= 8'h00;
		14'h1217:	ff_dbi <= 8'h00;
		14'h1218:	ff_dbi <= 8'h00;
		14'h1219:	ff_dbi <= 8'h00;
		14'h121a:	ff_dbi <= 8'h00;
		14'h121b:	ff_dbi <= 8'h00;
		14'h121c:	ff_dbi <= 8'h00;
		14'h121d:	ff_dbi <= 8'h00;
		14'h121e:	ff_dbi <= 8'h00;
		14'h121f:	ff_dbi <= 8'h00;
		14'h1220:	ff_dbi <= 8'h00;
		14'h1221:	ff_dbi <= 8'h00;
		14'h1222:	ff_dbi <= 8'h00;
		14'h1223:	ff_dbi <= 8'h00;
		14'h1224:	ff_dbi <= 8'h00;
		14'h1225:	ff_dbi <= 8'h00;
		14'h1226:	ff_dbi <= 8'h00;
		14'h1227:	ff_dbi <= 8'h00;
		14'h1228:	ff_dbi <= 8'h00;
		14'h1229:	ff_dbi <= 8'h00;
		14'h122a:	ff_dbi <= 8'h00;
		14'h122b:	ff_dbi <= 8'h00;
		14'h122c:	ff_dbi <= 8'h00;
		14'h122d:	ff_dbi <= 8'h00;
		14'h122e:	ff_dbi <= 8'h00;
		14'h122f:	ff_dbi <= 8'h00;
		14'h1230:	ff_dbi <= 8'h00;
		14'h1231:	ff_dbi <= 8'h00;
		14'h1232:	ff_dbi <= 8'h00;
		14'h1233:	ff_dbi <= 8'h00;
		14'h1234:	ff_dbi <= 8'h00;
		14'h1235:	ff_dbi <= 8'h00;
		14'h1236:	ff_dbi <= 8'h00;
		14'h1237:	ff_dbi <= 8'h00;
		14'h1238:	ff_dbi <= 8'h00;
		14'h1239:	ff_dbi <= 8'h00;
		14'h123a:	ff_dbi <= 8'h00;
		14'h123b:	ff_dbi <= 8'h00;
		14'h123c:	ff_dbi <= 8'h00;
		14'h123d:	ff_dbi <= 8'h00;
		14'h123e:	ff_dbi <= 8'h00;
		14'h123f:	ff_dbi <= 8'h00;
		14'h1240:	ff_dbi <= 8'h00;
		14'h1241:	ff_dbi <= 8'h00;
		14'h1242:	ff_dbi <= 8'h00;
		14'h1243:	ff_dbi <= 8'h00;
		14'h1244:	ff_dbi <= 8'h00;
		14'h1245:	ff_dbi <= 8'h00;
		14'h1246:	ff_dbi <= 8'h00;
		14'h1247:	ff_dbi <= 8'h00;
		14'h1248:	ff_dbi <= 8'h00;
		14'h1249:	ff_dbi <= 8'h00;
		14'h124a:	ff_dbi <= 8'h00;
		14'h124b:	ff_dbi <= 8'h00;
		14'h124c:	ff_dbi <= 8'h00;
		14'h124d:	ff_dbi <= 8'h00;
		14'h124e:	ff_dbi <= 8'h00;
		14'h124f:	ff_dbi <= 8'h00;
		14'h1250:	ff_dbi <= 8'h00;
		14'h1251:	ff_dbi <= 8'h00;
		14'h1252:	ff_dbi <= 8'h00;
		14'h1253:	ff_dbi <= 8'h00;
		14'h1254:	ff_dbi <= 8'h00;
		14'h1255:	ff_dbi <= 8'h00;
		14'h1256:	ff_dbi <= 8'h00;
		14'h1257:	ff_dbi <= 8'h00;
		14'h1258:	ff_dbi <= 8'h00;
		14'h1259:	ff_dbi <= 8'h00;
		14'h125a:	ff_dbi <= 8'h00;
		14'h125b:	ff_dbi <= 8'h00;
		14'h125c:	ff_dbi <= 8'h00;
		14'h125d:	ff_dbi <= 8'h00;
		14'h125e:	ff_dbi <= 8'h00;
		14'h125f:	ff_dbi <= 8'h00;
		14'h1260:	ff_dbi <= 8'h00;
		14'h1261:	ff_dbi <= 8'h00;
		14'h1262:	ff_dbi <= 8'h00;
		14'h1263:	ff_dbi <= 8'h00;
		14'h1264:	ff_dbi <= 8'h00;
		14'h1265:	ff_dbi <= 8'h00;
		14'h1266:	ff_dbi <= 8'h00;
		14'h1267:	ff_dbi <= 8'h00;
		14'h1268:	ff_dbi <= 8'h00;
		14'h1269:	ff_dbi <= 8'h00;
		14'h126a:	ff_dbi <= 8'h00;
		14'h126b:	ff_dbi <= 8'h00;
		14'h126c:	ff_dbi <= 8'h00;
		14'h126d:	ff_dbi <= 8'h00;
		14'h126e:	ff_dbi <= 8'h00;
		14'h126f:	ff_dbi <= 8'h00;
		14'h1270:	ff_dbi <= 8'h00;
		14'h1271:	ff_dbi <= 8'h00;
		14'h1272:	ff_dbi <= 8'h00;
		14'h1273:	ff_dbi <= 8'h00;
		14'h1274:	ff_dbi <= 8'h00;
		14'h1275:	ff_dbi <= 8'h00;
		14'h1276:	ff_dbi <= 8'h00;
		14'h1277:	ff_dbi <= 8'h00;
		14'h1278:	ff_dbi <= 8'h00;
		14'h1279:	ff_dbi <= 8'h00;
		14'h127a:	ff_dbi <= 8'h00;
		14'h127b:	ff_dbi <= 8'h00;
		14'h127c:	ff_dbi <= 8'h00;
		14'h127d:	ff_dbi <= 8'h00;
		14'h127e:	ff_dbi <= 8'h00;
		14'h127f:	ff_dbi <= 8'h00;
		14'h1280:	ff_dbi <= 8'h00;
		14'h1281:	ff_dbi <= 8'h00;
		14'h1282:	ff_dbi <= 8'h00;
		14'h1283:	ff_dbi <= 8'h00;
		14'h1284:	ff_dbi <= 8'h00;
		14'h1285:	ff_dbi <= 8'h00;
		14'h1286:	ff_dbi <= 8'h00;
		14'h1287:	ff_dbi <= 8'h00;
		14'h1288:	ff_dbi <= 8'h00;
		14'h1289:	ff_dbi <= 8'h00;
		14'h128a:	ff_dbi <= 8'h00;
		14'h128b:	ff_dbi <= 8'h00;
		14'h128c:	ff_dbi <= 8'h00;
		14'h128d:	ff_dbi <= 8'h00;
		14'h128e:	ff_dbi <= 8'h00;
		14'h128f:	ff_dbi <= 8'h00;
		14'h1290:	ff_dbi <= 8'h00;
		14'h1291:	ff_dbi <= 8'h00;
		14'h1292:	ff_dbi <= 8'h00;
		14'h1293:	ff_dbi <= 8'h00;
		14'h1294:	ff_dbi <= 8'h00;
		14'h1295:	ff_dbi <= 8'h00;
		14'h1296:	ff_dbi <= 8'h00;
		14'h1297:	ff_dbi <= 8'h00;
		14'h1298:	ff_dbi <= 8'h00;
		14'h1299:	ff_dbi <= 8'h00;
		14'h129a:	ff_dbi <= 8'h00;
		14'h129b:	ff_dbi <= 8'h00;
		14'h129c:	ff_dbi <= 8'h00;
		14'h129d:	ff_dbi <= 8'h00;
		14'h129e:	ff_dbi <= 8'h00;
		14'h129f:	ff_dbi <= 8'h00;
		14'h12a0:	ff_dbi <= 8'h00;
		14'h12a1:	ff_dbi <= 8'h00;
		14'h12a2:	ff_dbi <= 8'h00;
		14'h12a3:	ff_dbi <= 8'h00;
		14'h12a4:	ff_dbi <= 8'h00;
		14'h12a5:	ff_dbi <= 8'h00;
		14'h12a6:	ff_dbi <= 8'h00;
		14'h12a7:	ff_dbi <= 8'h00;
		14'h12a8:	ff_dbi <= 8'h00;
		14'h12a9:	ff_dbi <= 8'h00;
		14'h12aa:	ff_dbi <= 8'h00;
		14'h12ab:	ff_dbi <= 8'h00;
		14'h12ac:	ff_dbi <= 8'h00;
		14'h12ad:	ff_dbi <= 8'h00;
		14'h12ae:	ff_dbi <= 8'h00;
		14'h12af:	ff_dbi <= 8'h00;
		14'h12b0:	ff_dbi <= 8'h00;
		14'h12b1:	ff_dbi <= 8'h00;
		14'h12b2:	ff_dbi <= 8'h00;
		14'h12b3:	ff_dbi <= 8'h00;
		14'h12b4:	ff_dbi <= 8'h00;
		14'h12b5:	ff_dbi <= 8'h00;
		14'h12b6:	ff_dbi <= 8'h00;
		14'h12b7:	ff_dbi <= 8'h00;
		14'h12b8:	ff_dbi <= 8'h00;
		14'h12b9:	ff_dbi <= 8'h00;
		14'h12ba:	ff_dbi <= 8'h00;
		14'h12bb:	ff_dbi <= 8'h00;
		14'h12bc:	ff_dbi <= 8'h00;
		14'h12bd:	ff_dbi <= 8'h00;
		14'h12be:	ff_dbi <= 8'h00;
		14'h12bf:	ff_dbi <= 8'h00;
		14'h12c0:	ff_dbi <= 8'h00;
		14'h12c1:	ff_dbi <= 8'h00;
		14'h12c2:	ff_dbi <= 8'h00;
		14'h12c3:	ff_dbi <= 8'h00;
		14'h12c4:	ff_dbi <= 8'h00;
		14'h12c5:	ff_dbi <= 8'h00;
		14'h12c6:	ff_dbi <= 8'h00;
		14'h12c7:	ff_dbi <= 8'h00;
		14'h12c8:	ff_dbi <= 8'h00;
		14'h12c9:	ff_dbi <= 8'h00;
		14'h12ca:	ff_dbi <= 8'h00;
		14'h12cb:	ff_dbi <= 8'h00;
		14'h12cc:	ff_dbi <= 8'h00;
		14'h12cd:	ff_dbi <= 8'h00;
		14'h12ce:	ff_dbi <= 8'h00;
		14'h12cf:	ff_dbi <= 8'h00;
		14'h12d0:	ff_dbi <= 8'h00;
		14'h12d1:	ff_dbi <= 8'h00;
		14'h12d2:	ff_dbi <= 8'h00;
		14'h12d3:	ff_dbi <= 8'h00;
		14'h12d4:	ff_dbi <= 8'h00;
		14'h12d5:	ff_dbi <= 8'h00;
		14'h12d6:	ff_dbi <= 8'h00;
		14'h12d7:	ff_dbi <= 8'h00;
		14'h12d8:	ff_dbi <= 8'h00;
		14'h12d9:	ff_dbi <= 8'h00;
		14'h12da:	ff_dbi <= 8'h00;
		14'h12db:	ff_dbi <= 8'h00;
		14'h12dc:	ff_dbi <= 8'h00;
		14'h12dd:	ff_dbi <= 8'h00;
		14'h12de:	ff_dbi <= 8'h00;
		14'h12df:	ff_dbi <= 8'h00;
		14'h12e0:	ff_dbi <= 8'h00;
		14'h12e1:	ff_dbi <= 8'h00;
		14'h12e2:	ff_dbi <= 8'h00;
		14'h12e3:	ff_dbi <= 8'h00;
		14'h12e4:	ff_dbi <= 8'h00;
		14'h12e5:	ff_dbi <= 8'h00;
		14'h12e6:	ff_dbi <= 8'h00;
		14'h12e7:	ff_dbi <= 8'h00;
		14'h12e8:	ff_dbi <= 8'h00;
		14'h12e9:	ff_dbi <= 8'h00;
		14'h12ea:	ff_dbi <= 8'h00;
		14'h12eb:	ff_dbi <= 8'h00;
		14'h12ec:	ff_dbi <= 8'h00;
		14'h12ed:	ff_dbi <= 8'h00;
		14'h12ee:	ff_dbi <= 8'h00;
		14'h12ef:	ff_dbi <= 8'h00;
		14'h12f0:	ff_dbi <= 8'h00;
		14'h12f1:	ff_dbi <= 8'h00;
		14'h12f2:	ff_dbi <= 8'h00;
		14'h12f3:	ff_dbi <= 8'h00;
		14'h12f4:	ff_dbi <= 8'h00;
		14'h12f5:	ff_dbi <= 8'h00;
		14'h12f6:	ff_dbi <= 8'h00;
		14'h12f7:	ff_dbi <= 8'h00;
		14'h12f8:	ff_dbi <= 8'h00;
		14'h12f9:	ff_dbi <= 8'h00;
		14'h12fa:	ff_dbi <= 8'h00;
		14'h12fb:	ff_dbi <= 8'h00;
		14'h12fc:	ff_dbi <= 8'h00;
		14'h12fd:	ff_dbi <= 8'h00;
		14'h12fe:	ff_dbi <= 8'h00;
		14'h12ff:	ff_dbi <= 8'h00;
		14'h1300:	ff_dbi <= 8'h00;
		14'h1301:	ff_dbi <= 8'h00;
		14'h1302:	ff_dbi <= 8'h00;
		14'h1303:	ff_dbi <= 8'h00;
		14'h1304:	ff_dbi <= 8'h00;
		14'h1305:	ff_dbi <= 8'h00;
		14'h1306:	ff_dbi <= 8'h00;
		14'h1307:	ff_dbi <= 8'h00;
		14'h1308:	ff_dbi <= 8'h00;
		14'h1309:	ff_dbi <= 8'h00;
		14'h130a:	ff_dbi <= 8'h00;
		14'h130b:	ff_dbi <= 8'h00;
		14'h130c:	ff_dbi <= 8'h00;
		14'h130d:	ff_dbi <= 8'h00;
		14'h130e:	ff_dbi <= 8'h00;
		14'h130f:	ff_dbi <= 8'h00;
		14'h1310:	ff_dbi <= 8'h00;
		14'h1311:	ff_dbi <= 8'h00;
		14'h1312:	ff_dbi <= 8'h00;
		14'h1313:	ff_dbi <= 8'h00;
		14'h1314:	ff_dbi <= 8'h00;
		14'h1315:	ff_dbi <= 8'h00;
		14'h1316:	ff_dbi <= 8'h00;
		14'h1317:	ff_dbi <= 8'h00;
		14'h1318:	ff_dbi <= 8'h00;
		14'h1319:	ff_dbi <= 8'h00;
		14'h131a:	ff_dbi <= 8'h00;
		14'h131b:	ff_dbi <= 8'h00;
		14'h131c:	ff_dbi <= 8'h00;
		14'h131d:	ff_dbi <= 8'h00;
		14'h131e:	ff_dbi <= 8'h00;
		14'h131f:	ff_dbi <= 8'h00;
		14'h1320:	ff_dbi <= 8'h00;
		14'h1321:	ff_dbi <= 8'h00;
		14'h1322:	ff_dbi <= 8'h00;
		14'h1323:	ff_dbi <= 8'h00;
		14'h1324:	ff_dbi <= 8'h00;
		14'h1325:	ff_dbi <= 8'h00;
		14'h1326:	ff_dbi <= 8'h00;
		14'h1327:	ff_dbi <= 8'h00;
		14'h1328:	ff_dbi <= 8'h00;
		14'h1329:	ff_dbi <= 8'h00;
		14'h132a:	ff_dbi <= 8'h00;
		14'h132b:	ff_dbi <= 8'h00;
		14'h132c:	ff_dbi <= 8'h00;
		14'h132d:	ff_dbi <= 8'h00;
		14'h132e:	ff_dbi <= 8'h00;
		14'h132f:	ff_dbi <= 8'h00;
		14'h1330:	ff_dbi <= 8'h00;
		14'h1331:	ff_dbi <= 8'h00;
		14'h1332:	ff_dbi <= 8'h00;
		14'h1333:	ff_dbi <= 8'h00;
		14'h1334:	ff_dbi <= 8'h00;
		14'h1335:	ff_dbi <= 8'h00;
		14'h1336:	ff_dbi <= 8'h00;
		14'h1337:	ff_dbi <= 8'h00;
		14'h1338:	ff_dbi <= 8'h00;
		14'h1339:	ff_dbi <= 8'h00;
		14'h133a:	ff_dbi <= 8'h00;
		14'h133b:	ff_dbi <= 8'h00;
		14'h133c:	ff_dbi <= 8'h00;
		14'h133d:	ff_dbi <= 8'h00;
		14'h133e:	ff_dbi <= 8'h00;
		14'h133f:	ff_dbi <= 8'h00;
		14'h1340:	ff_dbi <= 8'h00;
		14'h1341:	ff_dbi <= 8'h00;
		14'h1342:	ff_dbi <= 8'h00;
		14'h1343:	ff_dbi <= 8'h00;
		14'h1344:	ff_dbi <= 8'h00;
		14'h1345:	ff_dbi <= 8'h00;
		14'h1346:	ff_dbi <= 8'h00;
		14'h1347:	ff_dbi <= 8'h00;
		14'h1348:	ff_dbi <= 8'h00;
		14'h1349:	ff_dbi <= 8'h00;
		14'h134a:	ff_dbi <= 8'h00;
		14'h134b:	ff_dbi <= 8'h00;
		14'h134c:	ff_dbi <= 8'h00;
		14'h134d:	ff_dbi <= 8'h00;
		14'h134e:	ff_dbi <= 8'h00;
		14'h134f:	ff_dbi <= 8'h00;
		14'h1350:	ff_dbi <= 8'h00;
		14'h1351:	ff_dbi <= 8'h00;
		14'h1352:	ff_dbi <= 8'h00;
		14'h1353:	ff_dbi <= 8'h00;
		14'h1354:	ff_dbi <= 8'h00;
		14'h1355:	ff_dbi <= 8'h00;
		14'h1356:	ff_dbi <= 8'h00;
		14'h1357:	ff_dbi <= 8'h00;
		14'h1358:	ff_dbi <= 8'h00;
		14'h1359:	ff_dbi <= 8'h00;
		14'h135a:	ff_dbi <= 8'h00;
		14'h135b:	ff_dbi <= 8'h00;
		14'h135c:	ff_dbi <= 8'h00;
		14'h135d:	ff_dbi <= 8'h00;
		14'h135e:	ff_dbi <= 8'h00;
		14'h135f:	ff_dbi <= 8'h00;
		14'h1360:	ff_dbi <= 8'h00;
		14'h1361:	ff_dbi <= 8'h00;
		14'h1362:	ff_dbi <= 8'h00;
		14'h1363:	ff_dbi <= 8'h00;
		14'h1364:	ff_dbi <= 8'h00;
		14'h1365:	ff_dbi <= 8'h00;
		14'h1366:	ff_dbi <= 8'h00;
		14'h1367:	ff_dbi <= 8'h00;
		14'h1368:	ff_dbi <= 8'h00;
		14'h1369:	ff_dbi <= 8'h00;
		14'h136a:	ff_dbi <= 8'h00;
		14'h136b:	ff_dbi <= 8'h00;
		14'h136c:	ff_dbi <= 8'h00;
		14'h136d:	ff_dbi <= 8'h00;
		14'h136e:	ff_dbi <= 8'h00;
		14'h136f:	ff_dbi <= 8'h00;
		14'h1370:	ff_dbi <= 8'h00;
		14'h1371:	ff_dbi <= 8'h00;
		14'h1372:	ff_dbi <= 8'h00;
		14'h1373:	ff_dbi <= 8'h00;
		14'h1374:	ff_dbi <= 8'h00;
		14'h1375:	ff_dbi <= 8'h00;
		14'h1376:	ff_dbi <= 8'h00;
		14'h1377:	ff_dbi <= 8'h00;
		14'h1378:	ff_dbi <= 8'h00;
		14'h1379:	ff_dbi <= 8'h00;
		14'h137a:	ff_dbi <= 8'h00;
		14'h137b:	ff_dbi <= 8'h00;
		14'h137c:	ff_dbi <= 8'h00;
		14'h137d:	ff_dbi <= 8'h00;
		14'h137e:	ff_dbi <= 8'h00;
		14'h137f:	ff_dbi <= 8'h00;
		14'h1380:	ff_dbi <= 8'h00;
		14'h1381:	ff_dbi <= 8'h00;
		14'h1382:	ff_dbi <= 8'h00;
		14'h1383:	ff_dbi <= 8'h00;
		14'h1384:	ff_dbi <= 8'h00;
		14'h1385:	ff_dbi <= 8'h00;
		14'h1386:	ff_dbi <= 8'h00;
		14'h1387:	ff_dbi <= 8'h00;
		14'h1388:	ff_dbi <= 8'h00;
		14'h1389:	ff_dbi <= 8'h00;
		14'h138a:	ff_dbi <= 8'h00;
		14'h138b:	ff_dbi <= 8'h00;
		14'h138c:	ff_dbi <= 8'h00;
		14'h138d:	ff_dbi <= 8'h00;
		14'h138e:	ff_dbi <= 8'h00;
		14'h138f:	ff_dbi <= 8'h00;
		14'h1390:	ff_dbi <= 8'h00;
		14'h1391:	ff_dbi <= 8'h00;
		14'h1392:	ff_dbi <= 8'h00;
		14'h1393:	ff_dbi <= 8'h00;
		14'h1394:	ff_dbi <= 8'h00;
		14'h1395:	ff_dbi <= 8'h00;
		14'h1396:	ff_dbi <= 8'h00;
		14'h1397:	ff_dbi <= 8'h00;
		14'h1398:	ff_dbi <= 8'h00;
		14'h1399:	ff_dbi <= 8'h00;
		14'h139a:	ff_dbi <= 8'h00;
		14'h139b:	ff_dbi <= 8'h00;
		14'h139c:	ff_dbi <= 8'h00;
		14'h139d:	ff_dbi <= 8'h00;
		14'h139e:	ff_dbi <= 8'h00;
		14'h139f:	ff_dbi <= 8'h00;
		14'h13a0:	ff_dbi <= 8'h00;
		14'h13a1:	ff_dbi <= 8'h00;
		14'h13a2:	ff_dbi <= 8'h00;
		14'h13a3:	ff_dbi <= 8'h00;
		14'h13a4:	ff_dbi <= 8'h00;
		14'h13a5:	ff_dbi <= 8'h00;
		14'h13a6:	ff_dbi <= 8'h00;
		14'h13a7:	ff_dbi <= 8'h00;
		14'h13a8:	ff_dbi <= 8'h00;
		14'h13a9:	ff_dbi <= 8'h00;
		14'h13aa:	ff_dbi <= 8'h00;
		14'h13ab:	ff_dbi <= 8'h00;
		14'h13ac:	ff_dbi <= 8'h00;
		14'h13ad:	ff_dbi <= 8'h00;
		14'h13ae:	ff_dbi <= 8'h00;
		14'h13af:	ff_dbi <= 8'h00;
		14'h13b0:	ff_dbi <= 8'h00;
		14'h13b1:	ff_dbi <= 8'h00;
		14'h13b2:	ff_dbi <= 8'h00;
		14'h13b3:	ff_dbi <= 8'h00;
		14'h13b4:	ff_dbi <= 8'h00;
		14'h13b5:	ff_dbi <= 8'h00;
		14'h13b6:	ff_dbi <= 8'h00;
		14'h13b7:	ff_dbi <= 8'h00;
		14'h13b8:	ff_dbi <= 8'h00;
		14'h13b9:	ff_dbi <= 8'h00;
		14'h13ba:	ff_dbi <= 8'h00;
		14'h13bb:	ff_dbi <= 8'h00;
		14'h13bc:	ff_dbi <= 8'h00;
		14'h13bd:	ff_dbi <= 8'h00;
		14'h13be:	ff_dbi <= 8'h00;
		14'h13bf:	ff_dbi <= 8'h00;
		14'h13c0:	ff_dbi <= 8'h00;
		14'h13c1:	ff_dbi <= 8'h00;
		14'h13c2:	ff_dbi <= 8'h00;
		14'h13c3:	ff_dbi <= 8'h00;
		14'h13c4:	ff_dbi <= 8'h00;
		14'h13c5:	ff_dbi <= 8'h00;
		14'h13c6:	ff_dbi <= 8'h00;
		14'h13c7:	ff_dbi <= 8'h00;
		14'h13c8:	ff_dbi <= 8'h00;
		14'h13c9:	ff_dbi <= 8'h00;
		14'h13ca:	ff_dbi <= 8'h00;
		14'h13cb:	ff_dbi <= 8'h00;
		14'h13cc:	ff_dbi <= 8'h00;
		14'h13cd:	ff_dbi <= 8'h00;
		14'h13ce:	ff_dbi <= 8'h00;
		14'h13cf:	ff_dbi <= 8'h00;
		14'h13d0:	ff_dbi <= 8'h00;
		14'h13d1:	ff_dbi <= 8'h00;
		14'h13d2:	ff_dbi <= 8'h00;
		14'h13d3:	ff_dbi <= 8'h00;
		14'h13d4:	ff_dbi <= 8'h00;
		14'h13d5:	ff_dbi <= 8'h00;
		14'h13d6:	ff_dbi <= 8'h00;
		14'h13d7:	ff_dbi <= 8'h00;
		14'h13d8:	ff_dbi <= 8'h00;
		14'h13d9:	ff_dbi <= 8'h00;
		14'h13da:	ff_dbi <= 8'h00;
		14'h13db:	ff_dbi <= 8'h00;
		14'h13dc:	ff_dbi <= 8'h00;
		14'h13dd:	ff_dbi <= 8'h00;
		14'h13de:	ff_dbi <= 8'h00;
		14'h13df:	ff_dbi <= 8'h00;
		14'h13e0:	ff_dbi <= 8'h00;
		14'h13e1:	ff_dbi <= 8'h00;
		14'h13e2:	ff_dbi <= 8'h00;
		14'h13e3:	ff_dbi <= 8'h00;
		14'h13e4:	ff_dbi <= 8'h00;
		14'h13e5:	ff_dbi <= 8'h00;
		14'h13e6:	ff_dbi <= 8'h00;
		14'h13e7:	ff_dbi <= 8'h00;
		14'h13e8:	ff_dbi <= 8'h00;
		14'h13e9:	ff_dbi <= 8'h00;
		14'h13ea:	ff_dbi <= 8'h00;
		14'h13eb:	ff_dbi <= 8'h00;
		14'h13ec:	ff_dbi <= 8'h00;
		14'h13ed:	ff_dbi <= 8'h00;
		14'h13ee:	ff_dbi <= 8'h00;
		14'h13ef:	ff_dbi <= 8'h00;
		14'h13f0:	ff_dbi <= 8'h00;
		14'h13f1:	ff_dbi <= 8'h00;
		14'h13f2:	ff_dbi <= 8'h00;
		14'h13f3:	ff_dbi <= 8'h00;
		14'h13f4:	ff_dbi <= 8'h00;
		14'h13f5:	ff_dbi <= 8'h00;
		14'h13f6:	ff_dbi <= 8'h00;
		14'h13f7:	ff_dbi <= 8'h00;
		14'h13f8:	ff_dbi <= 8'h00;
		14'h13f9:	ff_dbi <= 8'h00;
		14'h13fa:	ff_dbi <= 8'h00;
		14'h13fb:	ff_dbi <= 8'h00;
		14'h13fc:	ff_dbi <= 8'h00;
		14'h13fd:	ff_dbi <= 8'h00;
		14'h13fe:	ff_dbi <= 8'h00;
		14'h13ff:	ff_dbi <= 8'h00;
		14'h1400:	ff_dbi <= 8'h00;
		14'h1401:	ff_dbi <= 8'h00;
		14'h1402:	ff_dbi <= 8'h00;
		14'h1403:	ff_dbi <= 8'h00;
		14'h1404:	ff_dbi <= 8'h00;
		14'h1405:	ff_dbi <= 8'h00;
		14'h1406:	ff_dbi <= 8'h00;
		14'h1407:	ff_dbi <= 8'h00;
		14'h1408:	ff_dbi <= 8'h00;
		14'h1409:	ff_dbi <= 8'h00;
		14'h140a:	ff_dbi <= 8'h00;
		14'h140b:	ff_dbi <= 8'h00;
		14'h140c:	ff_dbi <= 8'h00;
		14'h140d:	ff_dbi <= 8'h00;
		14'h140e:	ff_dbi <= 8'h00;
		14'h140f:	ff_dbi <= 8'h00;
		14'h1410:	ff_dbi <= 8'h00;
		14'h1411:	ff_dbi <= 8'h00;
		14'h1412:	ff_dbi <= 8'h00;
		14'h1413:	ff_dbi <= 8'h00;
		14'h1414:	ff_dbi <= 8'h00;
		14'h1415:	ff_dbi <= 8'h00;
		14'h1416:	ff_dbi <= 8'h00;
		14'h1417:	ff_dbi <= 8'h00;
		14'h1418:	ff_dbi <= 8'h00;
		14'h1419:	ff_dbi <= 8'h00;
		14'h141a:	ff_dbi <= 8'h00;
		14'h141b:	ff_dbi <= 8'h00;
		14'h141c:	ff_dbi <= 8'h00;
		14'h141d:	ff_dbi <= 8'h00;
		14'h141e:	ff_dbi <= 8'h00;
		14'h141f:	ff_dbi <= 8'h00;
		14'h1420:	ff_dbi <= 8'h00;
		14'h1421:	ff_dbi <= 8'h00;
		14'h1422:	ff_dbi <= 8'h00;
		14'h1423:	ff_dbi <= 8'h00;
		14'h1424:	ff_dbi <= 8'h00;
		14'h1425:	ff_dbi <= 8'h00;
		14'h1426:	ff_dbi <= 8'h00;
		14'h1427:	ff_dbi <= 8'h00;
		14'h1428:	ff_dbi <= 8'h00;
		14'h1429:	ff_dbi <= 8'h00;
		14'h142a:	ff_dbi <= 8'h00;
		14'h142b:	ff_dbi <= 8'h00;
		14'h142c:	ff_dbi <= 8'h00;
		14'h142d:	ff_dbi <= 8'h00;
		14'h142e:	ff_dbi <= 8'h00;
		14'h142f:	ff_dbi <= 8'h00;
		14'h1430:	ff_dbi <= 8'h00;
		14'h1431:	ff_dbi <= 8'h00;
		14'h1432:	ff_dbi <= 8'h00;
		14'h1433:	ff_dbi <= 8'h00;
		14'h1434:	ff_dbi <= 8'h00;
		14'h1435:	ff_dbi <= 8'h00;
		14'h1436:	ff_dbi <= 8'h00;
		14'h1437:	ff_dbi <= 8'h00;
		14'h1438:	ff_dbi <= 8'h00;
		14'h1439:	ff_dbi <= 8'h00;
		14'h143a:	ff_dbi <= 8'h00;
		14'h143b:	ff_dbi <= 8'h00;
		14'h143c:	ff_dbi <= 8'h00;
		14'h143d:	ff_dbi <= 8'h00;
		14'h143e:	ff_dbi <= 8'h00;
		14'h143f:	ff_dbi <= 8'h00;
		14'h1440:	ff_dbi <= 8'h00;
		14'h1441:	ff_dbi <= 8'h00;
		14'h1442:	ff_dbi <= 8'h00;
		14'h1443:	ff_dbi <= 8'h00;
		14'h1444:	ff_dbi <= 8'h00;
		14'h1445:	ff_dbi <= 8'h00;
		14'h1446:	ff_dbi <= 8'h00;
		14'h1447:	ff_dbi <= 8'h00;
		14'h1448:	ff_dbi <= 8'h00;
		14'h1449:	ff_dbi <= 8'h00;
		14'h144a:	ff_dbi <= 8'h00;
		14'h144b:	ff_dbi <= 8'h00;
		14'h144c:	ff_dbi <= 8'h00;
		14'h144d:	ff_dbi <= 8'h00;
		14'h144e:	ff_dbi <= 8'h00;
		14'h144f:	ff_dbi <= 8'h00;
		14'h1450:	ff_dbi <= 8'h00;
		14'h1451:	ff_dbi <= 8'h00;
		14'h1452:	ff_dbi <= 8'h00;
		14'h1453:	ff_dbi <= 8'h00;
		14'h1454:	ff_dbi <= 8'h00;
		14'h1455:	ff_dbi <= 8'h00;
		14'h1456:	ff_dbi <= 8'h00;
		14'h1457:	ff_dbi <= 8'h00;
		14'h1458:	ff_dbi <= 8'h00;
		14'h1459:	ff_dbi <= 8'h00;
		14'h145a:	ff_dbi <= 8'h00;
		14'h145b:	ff_dbi <= 8'h00;
		14'h145c:	ff_dbi <= 8'h00;
		14'h145d:	ff_dbi <= 8'h00;
		14'h145e:	ff_dbi <= 8'h00;
		14'h145f:	ff_dbi <= 8'h00;
		14'h1460:	ff_dbi <= 8'h00;
		14'h1461:	ff_dbi <= 8'h00;
		14'h1462:	ff_dbi <= 8'h00;
		14'h1463:	ff_dbi <= 8'h00;
		14'h1464:	ff_dbi <= 8'h00;
		14'h1465:	ff_dbi <= 8'h00;
		14'h1466:	ff_dbi <= 8'h00;
		14'h1467:	ff_dbi <= 8'h00;
		14'h1468:	ff_dbi <= 8'h00;
		14'h1469:	ff_dbi <= 8'h00;
		14'h146a:	ff_dbi <= 8'h00;
		14'h146b:	ff_dbi <= 8'h00;
		14'h146c:	ff_dbi <= 8'h00;
		14'h146d:	ff_dbi <= 8'h00;
		14'h146e:	ff_dbi <= 8'h00;
		14'h146f:	ff_dbi <= 8'h00;
		14'h1470:	ff_dbi <= 8'h00;
		14'h1471:	ff_dbi <= 8'h00;
		14'h1472:	ff_dbi <= 8'h00;
		14'h1473:	ff_dbi <= 8'h00;
		14'h1474:	ff_dbi <= 8'h00;
		14'h1475:	ff_dbi <= 8'h00;
		14'h1476:	ff_dbi <= 8'h00;
		14'h1477:	ff_dbi <= 8'h00;
		14'h1478:	ff_dbi <= 8'h00;
		14'h1479:	ff_dbi <= 8'h00;
		14'h147a:	ff_dbi <= 8'h00;
		14'h147b:	ff_dbi <= 8'h00;
		14'h147c:	ff_dbi <= 8'h00;
		14'h147d:	ff_dbi <= 8'h00;
		14'h147e:	ff_dbi <= 8'h00;
		14'h147f:	ff_dbi <= 8'h00;
		14'h1480:	ff_dbi <= 8'h00;
		14'h1481:	ff_dbi <= 8'h00;
		14'h1482:	ff_dbi <= 8'h00;
		14'h1483:	ff_dbi <= 8'h00;
		14'h1484:	ff_dbi <= 8'h00;
		14'h1485:	ff_dbi <= 8'h00;
		14'h1486:	ff_dbi <= 8'h00;
		14'h1487:	ff_dbi <= 8'h00;
		14'h1488:	ff_dbi <= 8'h00;
		14'h1489:	ff_dbi <= 8'h00;
		14'h148a:	ff_dbi <= 8'h00;
		14'h148b:	ff_dbi <= 8'h00;
		14'h148c:	ff_dbi <= 8'h00;
		14'h148d:	ff_dbi <= 8'h00;
		14'h148e:	ff_dbi <= 8'h00;
		14'h148f:	ff_dbi <= 8'h00;
		14'h1490:	ff_dbi <= 8'h00;
		14'h1491:	ff_dbi <= 8'h00;
		14'h1492:	ff_dbi <= 8'h00;
		14'h1493:	ff_dbi <= 8'h00;
		14'h1494:	ff_dbi <= 8'h00;
		14'h1495:	ff_dbi <= 8'h00;
		14'h1496:	ff_dbi <= 8'h00;
		14'h1497:	ff_dbi <= 8'h00;
		14'h1498:	ff_dbi <= 8'h00;
		14'h1499:	ff_dbi <= 8'h00;
		14'h149a:	ff_dbi <= 8'h00;
		14'h149b:	ff_dbi <= 8'h00;
		14'h149c:	ff_dbi <= 8'h00;
		14'h149d:	ff_dbi <= 8'h00;
		14'h149e:	ff_dbi <= 8'h00;
		14'h149f:	ff_dbi <= 8'h00;
		14'h14a0:	ff_dbi <= 8'h00;
		14'h14a1:	ff_dbi <= 8'h00;
		14'h14a2:	ff_dbi <= 8'h00;
		14'h14a3:	ff_dbi <= 8'h00;
		14'h14a4:	ff_dbi <= 8'h00;
		14'h14a5:	ff_dbi <= 8'h00;
		14'h14a6:	ff_dbi <= 8'h00;
		14'h14a7:	ff_dbi <= 8'h00;
		14'h14a8:	ff_dbi <= 8'h00;
		14'h14a9:	ff_dbi <= 8'h00;
		14'h14aa:	ff_dbi <= 8'h00;
		14'h14ab:	ff_dbi <= 8'h00;
		14'h14ac:	ff_dbi <= 8'h00;
		14'h14ad:	ff_dbi <= 8'h00;
		14'h14ae:	ff_dbi <= 8'h00;
		14'h14af:	ff_dbi <= 8'h00;
		14'h14b0:	ff_dbi <= 8'h00;
		14'h14b1:	ff_dbi <= 8'h00;
		14'h14b2:	ff_dbi <= 8'h00;
		14'h14b3:	ff_dbi <= 8'h00;
		14'h14b4:	ff_dbi <= 8'h00;
		14'h14b5:	ff_dbi <= 8'h00;
		14'h14b6:	ff_dbi <= 8'h00;
		14'h14b7:	ff_dbi <= 8'h00;
		14'h14b8:	ff_dbi <= 8'h00;
		14'h14b9:	ff_dbi <= 8'h00;
		14'h14ba:	ff_dbi <= 8'h00;
		14'h14bb:	ff_dbi <= 8'h00;
		14'h14bc:	ff_dbi <= 8'h00;
		14'h14bd:	ff_dbi <= 8'h00;
		14'h14be:	ff_dbi <= 8'h00;
		14'h14bf:	ff_dbi <= 8'h00;
		14'h14c0:	ff_dbi <= 8'h00;
		14'h14c1:	ff_dbi <= 8'h00;
		14'h14c2:	ff_dbi <= 8'h00;
		14'h14c3:	ff_dbi <= 8'h00;
		14'h14c4:	ff_dbi <= 8'h00;
		14'h14c5:	ff_dbi <= 8'h00;
		14'h14c6:	ff_dbi <= 8'h00;
		14'h14c7:	ff_dbi <= 8'h00;
		14'h14c8:	ff_dbi <= 8'h00;
		14'h14c9:	ff_dbi <= 8'h00;
		14'h14ca:	ff_dbi <= 8'h00;
		14'h14cb:	ff_dbi <= 8'h00;
		14'h14cc:	ff_dbi <= 8'h00;
		14'h14cd:	ff_dbi <= 8'h00;
		14'h14ce:	ff_dbi <= 8'h00;
		14'h14cf:	ff_dbi <= 8'h00;
		14'h14d0:	ff_dbi <= 8'h00;
		14'h14d1:	ff_dbi <= 8'h00;
		14'h14d2:	ff_dbi <= 8'h00;
		14'h14d3:	ff_dbi <= 8'h00;
		14'h14d4:	ff_dbi <= 8'h00;
		14'h14d5:	ff_dbi <= 8'h00;
		14'h14d6:	ff_dbi <= 8'h00;
		14'h14d7:	ff_dbi <= 8'h00;
		14'h14d8:	ff_dbi <= 8'h00;
		14'h14d9:	ff_dbi <= 8'h00;
		14'h14da:	ff_dbi <= 8'h00;
		14'h14db:	ff_dbi <= 8'h00;
		14'h14dc:	ff_dbi <= 8'h00;
		14'h14dd:	ff_dbi <= 8'h00;
		14'h14de:	ff_dbi <= 8'h00;
		14'h14df:	ff_dbi <= 8'h00;
		14'h14e0:	ff_dbi <= 8'h00;
		14'h14e1:	ff_dbi <= 8'h00;
		14'h14e2:	ff_dbi <= 8'h00;
		14'h14e3:	ff_dbi <= 8'h00;
		14'h14e4:	ff_dbi <= 8'h00;
		14'h14e5:	ff_dbi <= 8'h00;
		14'h14e6:	ff_dbi <= 8'h00;
		14'h14e7:	ff_dbi <= 8'h00;
		14'h14e8:	ff_dbi <= 8'h00;
		14'h14e9:	ff_dbi <= 8'h00;
		14'h14ea:	ff_dbi <= 8'h00;
		14'h14eb:	ff_dbi <= 8'h00;
		14'h14ec:	ff_dbi <= 8'h00;
		14'h14ed:	ff_dbi <= 8'h00;
		14'h14ee:	ff_dbi <= 8'h00;
		14'h14ef:	ff_dbi <= 8'h00;
		14'h14f0:	ff_dbi <= 8'h00;
		14'h14f1:	ff_dbi <= 8'h00;
		14'h14f2:	ff_dbi <= 8'h00;
		14'h14f3:	ff_dbi <= 8'h00;
		14'h14f4:	ff_dbi <= 8'h00;
		14'h14f5:	ff_dbi <= 8'h00;
		14'h14f6:	ff_dbi <= 8'h00;
		14'h14f7:	ff_dbi <= 8'h00;
		14'h14f8:	ff_dbi <= 8'h00;
		14'h14f9:	ff_dbi <= 8'h00;
		14'h14fa:	ff_dbi <= 8'h00;
		14'h14fb:	ff_dbi <= 8'h00;
		14'h14fc:	ff_dbi <= 8'h00;
		14'h14fd:	ff_dbi <= 8'h00;
		14'h14fe:	ff_dbi <= 8'h00;
		14'h14ff:	ff_dbi <= 8'h00;
		14'h1500:	ff_dbi <= 8'h00;
		14'h1501:	ff_dbi <= 8'h00;
		14'h1502:	ff_dbi <= 8'h00;
		14'h1503:	ff_dbi <= 8'h00;
		14'h1504:	ff_dbi <= 8'h00;
		14'h1505:	ff_dbi <= 8'h00;
		14'h1506:	ff_dbi <= 8'h00;
		14'h1507:	ff_dbi <= 8'h00;
		14'h1508:	ff_dbi <= 8'h00;
		14'h1509:	ff_dbi <= 8'h00;
		14'h150a:	ff_dbi <= 8'h00;
		14'h150b:	ff_dbi <= 8'h00;
		14'h150c:	ff_dbi <= 8'h00;
		14'h150d:	ff_dbi <= 8'h00;
		14'h150e:	ff_dbi <= 8'h00;
		14'h150f:	ff_dbi <= 8'h00;
		14'h1510:	ff_dbi <= 8'h00;
		14'h1511:	ff_dbi <= 8'h00;
		14'h1512:	ff_dbi <= 8'h00;
		14'h1513:	ff_dbi <= 8'h00;
		14'h1514:	ff_dbi <= 8'h00;
		14'h1515:	ff_dbi <= 8'h00;
		14'h1516:	ff_dbi <= 8'h00;
		14'h1517:	ff_dbi <= 8'h00;
		14'h1518:	ff_dbi <= 8'h00;
		14'h1519:	ff_dbi <= 8'h00;
		14'h151a:	ff_dbi <= 8'h00;
		14'h151b:	ff_dbi <= 8'h00;
		14'h151c:	ff_dbi <= 8'h00;
		14'h151d:	ff_dbi <= 8'h00;
		14'h151e:	ff_dbi <= 8'h00;
		14'h151f:	ff_dbi <= 8'h00;
		14'h1520:	ff_dbi <= 8'h00;
		14'h1521:	ff_dbi <= 8'h00;
		14'h1522:	ff_dbi <= 8'h00;
		14'h1523:	ff_dbi <= 8'h00;
		14'h1524:	ff_dbi <= 8'h00;
		14'h1525:	ff_dbi <= 8'h00;
		14'h1526:	ff_dbi <= 8'h00;
		14'h1527:	ff_dbi <= 8'h00;
		14'h1528:	ff_dbi <= 8'h00;
		14'h1529:	ff_dbi <= 8'h00;
		14'h152a:	ff_dbi <= 8'h00;
		14'h152b:	ff_dbi <= 8'h00;
		14'h152c:	ff_dbi <= 8'h00;
		14'h152d:	ff_dbi <= 8'h00;
		14'h152e:	ff_dbi <= 8'h00;
		14'h152f:	ff_dbi <= 8'h00;
		14'h1530:	ff_dbi <= 8'h00;
		14'h1531:	ff_dbi <= 8'h00;
		14'h1532:	ff_dbi <= 8'h00;
		14'h1533:	ff_dbi <= 8'h00;
		14'h1534:	ff_dbi <= 8'h00;
		14'h1535:	ff_dbi <= 8'h00;
		14'h1536:	ff_dbi <= 8'h00;
		14'h1537:	ff_dbi <= 8'h00;
		14'h1538:	ff_dbi <= 8'h00;
		14'h1539:	ff_dbi <= 8'h00;
		14'h153a:	ff_dbi <= 8'h00;
		14'h153b:	ff_dbi <= 8'h00;
		14'h153c:	ff_dbi <= 8'h00;
		14'h153d:	ff_dbi <= 8'h00;
		14'h153e:	ff_dbi <= 8'h00;
		14'h153f:	ff_dbi <= 8'h00;
		14'h1540:	ff_dbi <= 8'h00;
		14'h1541:	ff_dbi <= 8'h00;
		14'h1542:	ff_dbi <= 8'h00;
		14'h1543:	ff_dbi <= 8'h00;
		14'h1544:	ff_dbi <= 8'h00;
		14'h1545:	ff_dbi <= 8'h00;
		14'h1546:	ff_dbi <= 8'h00;
		14'h1547:	ff_dbi <= 8'h00;
		14'h1548:	ff_dbi <= 8'h00;
		14'h1549:	ff_dbi <= 8'h00;
		14'h154a:	ff_dbi <= 8'h00;
		14'h154b:	ff_dbi <= 8'h00;
		14'h154c:	ff_dbi <= 8'h00;
		14'h154d:	ff_dbi <= 8'h00;
		14'h154e:	ff_dbi <= 8'h00;
		14'h154f:	ff_dbi <= 8'h00;
		14'h1550:	ff_dbi <= 8'h00;
		14'h1551:	ff_dbi <= 8'h00;
		14'h1552:	ff_dbi <= 8'h00;
		14'h1553:	ff_dbi <= 8'h00;
		14'h1554:	ff_dbi <= 8'h00;
		14'h1555:	ff_dbi <= 8'h00;
		14'h1556:	ff_dbi <= 8'h00;
		14'h1557:	ff_dbi <= 8'h00;
		14'h1558:	ff_dbi <= 8'h00;
		14'h1559:	ff_dbi <= 8'h00;
		14'h155a:	ff_dbi <= 8'h00;
		14'h155b:	ff_dbi <= 8'h00;
		14'h155c:	ff_dbi <= 8'h00;
		14'h155d:	ff_dbi <= 8'h00;
		14'h155e:	ff_dbi <= 8'h00;
		14'h155f:	ff_dbi <= 8'h00;
		14'h1560:	ff_dbi <= 8'h00;
		14'h1561:	ff_dbi <= 8'h00;
		14'h1562:	ff_dbi <= 8'h00;
		14'h1563:	ff_dbi <= 8'h00;
		14'h1564:	ff_dbi <= 8'h00;
		14'h1565:	ff_dbi <= 8'h00;
		14'h1566:	ff_dbi <= 8'h00;
		14'h1567:	ff_dbi <= 8'h00;
		14'h1568:	ff_dbi <= 8'h00;
		14'h1569:	ff_dbi <= 8'h00;
		14'h156a:	ff_dbi <= 8'h00;
		14'h156b:	ff_dbi <= 8'h00;
		14'h156c:	ff_dbi <= 8'h00;
		14'h156d:	ff_dbi <= 8'h00;
		14'h156e:	ff_dbi <= 8'h00;
		14'h156f:	ff_dbi <= 8'h00;
		14'h1570:	ff_dbi <= 8'h00;
		14'h1571:	ff_dbi <= 8'h00;
		14'h1572:	ff_dbi <= 8'h00;
		14'h1573:	ff_dbi <= 8'h00;
		14'h1574:	ff_dbi <= 8'h00;
		14'h1575:	ff_dbi <= 8'h00;
		14'h1576:	ff_dbi <= 8'h00;
		14'h1577:	ff_dbi <= 8'h00;
		14'h1578:	ff_dbi <= 8'h00;
		14'h1579:	ff_dbi <= 8'h00;
		14'h157a:	ff_dbi <= 8'h00;
		14'h157b:	ff_dbi <= 8'h00;
		14'h157c:	ff_dbi <= 8'h00;
		14'h157d:	ff_dbi <= 8'h00;
		14'h157e:	ff_dbi <= 8'h00;
		14'h157f:	ff_dbi <= 8'h00;
		14'h1580:	ff_dbi <= 8'h00;
		14'h1581:	ff_dbi <= 8'h00;
		14'h1582:	ff_dbi <= 8'h00;
		14'h1583:	ff_dbi <= 8'h00;
		14'h1584:	ff_dbi <= 8'h00;
		14'h1585:	ff_dbi <= 8'h00;
		14'h1586:	ff_dbi <= 8'h00;
		14'h1587:	ff_dbi <= 8'h00;
		14'h1588:	ff_dbi <= 8'h00;
		14'h1589:	ff_dbi <= 8'h00;
		14'h158a:	ff_dbi <= 8'h00;
		14'h158b:	ff_dbi <= 8'h00;
		14'h158c:	ff_dbi <= 8'h00;
		14'h158d:	ff_dbi <= 8'h00;
		14'h158e:	ff_dbi <= 8'h00;
		14'h158f:	ff_dbi <= 8'h00;
		14'h1590:	ff_dbi <= 8'h00;
		14'h1591:	ff_dbi <= 8'h00;
		14'h1592:	ff_dbi <= 8'h00;
		14'h1593:	ff_dbi <= 8'h00;
		14'h1594:	ff_dbi <= 8'h00;
		14'h1595:	ff_dbi <= 8'h00;
		14'h1596:	ff_dbi <= 8'h00;
		14'h1597:	ff_dbi <= 8'h00;
		14'h1598:	ff_dbi <= 8'h00;
		14'h1599:	ff_dbi <= 8'h00;
		14'h159a:	ff_dbi <= 8'h00;
		14'h159b:	ff_dbi <= 8'h00;
		14'h159c:	ff_dbi <= 8'h00;
		14'h159d:	ff_dbi <= 8'h00;
		14'h159e:	ff_dbi <= 8'h00;
		14'h159f:	ff_dbi <= 8'h00;
		14'h15a0:	ff_dbi <= 8'h00;
		14'h15a1:	ff_dbi <= 8'h00;
		14'h15a2:	ff_dbi <= 8'h00;
		14'h15a3:	ff_dbi <= 8'h00;
		14'h15a4:	ff_dbi <= 8'h00;
		14'h15a5:	ff_dbi <= 8'h00;
		14'h15a6:	ff_dbi <= 8'h00;
		14'h15a7:	ff_dbi <= 8'h00;
		14'h15a8:	ff_dbi <= 8'h00;
		14'h15a9:	ff_dbi <= 8'h00;
		14'h15aa:	ff_dbi <= 8'h00;
		14'h15ab:	ff_dbi <= 8'h00;
		14'h15ac:	ff_dbi <= 8'h00;
		14'h15ad:	ff_dbi <= 8'h00;
		14'h15ae:	ff_dbi <= 8'h00;
		14'h15af:	ff_dbi <= 8'h00;
		14'h15b0:	ff_dbi <= 8'h00;
		14'h15b1:	ff_dbi <= 8'h00;
		14'h15b2:	ff_dbi <= 8'h00;
		14'h15b3:	ff_dbi <= 8'h00;
		14'h15b4:	ff_dbi <= 8'h00;
		14'h15b5:	ff_dbi <= 8'h00;
		14'h15b6:	ff_dbi <= 8'h00;
		14'h15b7:	ff_dbi <= 8'h00;
		14'h15b8:	ff_dbi <= 8'h00;
		14'h15b9:	ff_dbi <= 8'h00;
		14'h15ba:	ff_dbi <= 8'h00;
		14'h15bb:	ff_dbi <= 8'h00;
		14'h15bc:	ff_dbi <= 8'h00;
		14'h15bd:	ff_dbi <= 8'h00;
		14'h15be:	ff_dbi <= 8'h00;
		14'h15bf:	ff_dbi <= 8'h00;
		14'h15c0:	ff_dbi <= 8'h00;
		14'h15c1:	ff_dbi <= 8'h00;
		14'h15c2:	ff_dbi <= 8'h00;
		14'h15c3:	ff_dbi <= 8'h00;
		14'h15c4:	ff_dbi <= 8'h00;
		14'h15c5:	ff_dbi <= 8'h00;
		14'h15c6:	ff_dbi <= 8'h00;
		14'h15c7:	ff_dbi <= 8'h00;
		14'h15c8:	ff_dbi <= 8'h00;
		14'h15c9:	ff_dbi <= 8'h00;
		14'h15ca:	ff_dbi <= 8'h00;
		14'h15cb:	ff_dbi <= 8'h00;
		14'h15cc:	ff_dbi <= 8'h00;
		14'h15cd:	ff_dbi <= 8'h00;
		14'h15ce:	ff_dbi <= 8'h00;
		14'h15cf:	ff_dbi <= 8'h00;
		14'h15d0:	ff_dbi <= 8'h00;
		14'h15d1:	ff_dbi <= 8'h00;
		14'h15d2:	ff_dbi <= 8'h00;
		14'h15d3:	ff_dbi <= 8'h00;
		14'h15d4:	ff_dbi <= 8'h00;
		14'h15d5:	ff_dbi <= 8'h00;
		14'h15d6:	ff_dbi <= 8'h00;
		14'h15d7:	ff_dbi <= 8'h00;
		14'h15d8:	ff_dbi <= 8'h00;
		14'h15d9:	ff_dbi <= 8'h00;
		14'h15da:	ff_dbi <= 8'h00;
		14'h15db:	ff_dbi <= 8'h00;
		14'h15dc:	ff_dbi <= 8'h00;
		14'h15dd:	ff_dbi <= 8'h00;
		14'h15de:	ff_dbi <= 8'h00;
		14'h15df:	ff_dbi <= 8'h00;
		14'h15e0:	ff_dbi <= 8'h00;
		14'h15e1:	ff_dbi <= 8'h00;
		14'h15e2:	ff_dbi <= 8'h00;
		14'h15e3:	ff_dbi <= 8'h00;
		14'h15e4:	ff_dbi <= 8'h00;
		14'h15e5:	ff_dbi <= 8'h00;
		14'h15e6:	ff_dbi <= 8'h00;
		14'h15e7:	ff_dbi <= 8'h00;
		14'h15e8:	ff_dbi <= 8'h00;
		14'h15e9:	ff_dbi <= 8'h00;
		14'h15ea:	ff_dbi <= 8'h00;
		14'h15eb:	ff_dbi <= 8'h00;
		14'h15ec:	ff_dbi <= 8'h00;
		14'h15ed:	ff_dbi <= 8'h00;
		14'h15ee:	ff_dbi <= 8'h00;
		14'h15ef:	ff_dbi <= 8'h00;
		14'h15f0:	ff_dbi <= 8'h00;
		14'h15f1:	ff_dbi <= 8'h00;
		14'h15f2:	ff_dbi <= 8'h00;
		14'h15f3:	ff_dbi <= 8'h00;
		14'h15f4:	ff_dbi <= 8'h00;
		14'h15f5:	ff_dbi <= 8'h00;
		14'h15f6:	ff_dbi <= 8'h00;
		14'h15f7:	ff_dbi <= 8'h00;
		14'h15f8:	ff_dbi <= 8'h00;
		14'h15f9:	ff_dbi <= 8'h00;
		14'h15fa:	ff_dbi <= 8'h00;
		14'h15fb:	ff_dbi <= 8'h00;
		14'h15fc:	ff_dbi <= 8'h00;
		14'h15fd:	ff_dbi <= 8'h00;
		14'h15fe:	ff_dbi <= 8'h00;
		14'h15ff:	ff_dbi <= 8'h00;
		14'h1600:	ff_dbi <= 8'h00;
		14'h1601:	ff_dbi <= 8'h00;
		14'h1602:	ff_dbi <= 8'h00;
		14'h1603:	ff_dbi <= 8'h00;
		14'h1604:	ff_dbi <= 8'h00;
		14'h1605:	ff_dbi <= 8'h00;
		14'h1606:	ff_dbi <= 8'h00;
		14'h1607:	ff_dbi <= 8'h00;
		14'h1608:	ff_dbi <= 8'h00;
		14'h1609:	ff_dbi <= 8'h00;
		14'h160a:	ff_dbi <= 8'h00;
		14'h160b:	ff_dbi <= 8'h00;
		14'h160c:	ff_dbi <= 8'h00;
		14'h160d:	ff_dbi <= 8'h00;
		14'h160e:	ff_dbi <= 8'h00;
		14'h160f:	ff_dbi <= 8'h00;
		14'h1610:	ff_dbi <= 8'h00;
		14'h1611:	ff_dbi <= 8'h00;
		14'h1612:	ff_dbi <= 8'h00;
		14'h1613:	ff_dbi <= 8'h00;
		14'h1614:	ff_dbi <= 8'h00;
		14'h1615:	ff_dbi <= 8'h00;
		14'h1616:	ff_dbi <= 8'h00;
		14'h1617:	ff_dbi <= 8'h00;
		14'h1618:	ff_dbi <= 8'h00;
		14'h1619:	ff_dbi <= 8'h00;
		14'h161a:	ff_dbi <= 8'h00;
		14'h161b:	ff_dbi <= 8'h00;
		14'h161c:	ff_dbi <= 8'h00;
		14'h161d:	ff_dbi <= 8'h00;
		14'h161e:	ff_dbi <= 8'h00;
		14'h161f:	ff_dbi <= 8'h00;
		14'h1620:	ff_dbi <= 8'h00;
		14'h1621:	ff_dbi <= 8'h00;
		14'h1622:	ff_dbi <= 8'h00;
		14'h1623:	ff_dbi <= 8'h00;
		14'h1624:	ff_dbi <= 8'h00;
		14'h1625:	ff_dbi <= 8'h00;
		14'h1626:	ff_dbi <= 8'h00;
		14'h1627:	ff_dbi <= 8'h00;
		14'h1628:	ff_dbi <= 8'h00;
		14'h1629:	ff_dbi <= 8'h00;
		14'h162a:	ff_dbi <= 8'h00;
		14'h162b:	ff_dbi <= 8'h00;
		14'h162c:	ff_dbi <= 8'h00;
		14'h162d:	ff_dbi <= 8'h00;
		14'h162e:	ff_dbi <= 8'h00;
		14'h162f:	ff_dbi <= 8'h00;
		14'h1630:	ff_dbi <= 8'h00;
		14'h1631:	ff_dbi <= 8'h00;
		14'h1632:	ff_dbi <= 8'h00;
		14'h1633:	ff_dbi <= 8'h00;
		14'h1634:	ff_dbi <= 8'h00;
		14'h1635:	ff_dbi <= 8'h00;
		14'h1636:	ff_dbi <= 8'h00;
		14'h1637:	ff_dbi <= 8'h00;
		14'h1638:	ff_dbi <= 8'h00;
		14'h1639:	ff_dbi <= 8'h00;
		14'h163a:	ff_dbi <= 8'h00;
		14'h163b:	ff_dbi <= 8'h00;
		14'h163c:	ff_dbi <= 8'h00;
		14'h163d:	ff_dbi <= 8'h00;
		14'h163e:	ff_dbi <= 8'h00;
		14'h163f:	ff_dbi <= 8'h00;
		14'h1640:	ff_dbi <= 8'h00;
		14'h1641:	ff_dbi <= 8'h00;
		14'h1642:	ff_dbi <= 8'h00;
		14'h1643:	ff_dbi <= 8'h00;
		14'h1644:	ff_dbi <= 8'h00;
		14'h1645:	ff_dbi <= 8'h00;
		14'h1646:	ff_dbi <= 8'h00;
		14'h1647:	ff_dbi <= 8'h00;
		14'h1648:	ff_dbi <= 8'h00;
		14'h1649:	ff_dbi <= 8'h00;
		14'h164a:	ff_dbi <= 8'h00;
		14'h164b:	ff_dbi <= 8'h00;
		14'h164c:	ff_dbi <= 8'h00;
		14'h164d:	ff_dbi <= 8'h00;
		14'h164e:	ff_dbi <= 8'h00;
		14'h164f:	ff_dbi <= 8'h00;
		14'h1650:	ff_dbi <= 8'h00;
		14'h1651:	ff_dbi <= 8'h00;
		14'h1652:	ff_dbi <= 8'h00;
		14'h1653:	ff_dbi <= 8'h00;
		14'h1654:	ff_dbi <= 8'h00;
		14'h1655:	ff_dbi <= 8'h00;
		14'h1656:	ff_dbi <= 8'h00;
		14'h1657:	ff_dbi <= 8'h00;
		14'h1658:	ff_dbi <= 8'h00;
		14'h1659:	ff_dbi <= 8'h00;
		14'h165a:	ff_dbi <= 8'h00;
		14'h165b:	ff_dbi <= 8'h00;
		14'h165c:	ff_dbi <= 8'h00;
		14'h165d:	ff_dbi <= 8'h00;
		14'h165e:	ff_dbi <= 8'h00;
		14'h165f:	ff_dbi <= 8'h00;
		14'h1660:	ff_dbi <= 8'h00;
		14'h1661:	ff_dbi <= 8'h00;
		14'h1662:	ff_dbi <= 8'h00;
		14'h1663:	ff_dbi <= 8'h00;
		14'h1664:	ff_dbi <= 8'h00;
		14'h1665:	ff_dbi <= 8'h00;
		14'h1666:	ff_dbi <= 8'h00;
		14'h1667:	ff_dbi <= 8'h00;
		14'h1668:	ff_dbi <= 8'h00;
		14'h1669:	ff_dbi <= 8'h00;
		14'h166a:	ff_dbi <= 8'h00;
		14'h166b:	ff_dbi <= 8'h00;
		14'h166c:	ff_dbi <= 8'h00;
		14'h166d:	ff_dbi <= 8'h00;
		14'h166e:	ff_dbi <= 8'h00;
		14'h166f:	ff_dbi <= 8'h00;
		14'h1670:	ff_dbi <= 8'h00;
		14'h1671:	ff_dbi <= 8'h00;
		14'h1672:	ff_dbi <= 8'h00;
		14'h1673:	ff_dbi <= 8'h00;
		14'h1674:	ff_dbi <= 8'h00;
		14'h1675:	ff_dbi <= 8'h00;
		14'h1676:	ff_dbi <= 8'h00;
		14'h1677:	ff_dbi <= 8'h00;
		14'h1678:	ff_dbi <= 8'h00;
		14'h1679:	ff_dbi <= 8'h00;
		14'h167a:	ff_dbi <= 8'h00;
		14'h167b:	ff_dbi <= 8'h00;
		14'h167c:	ff_dbi <= 8'h00;
		14'h167d:	ff_dbi <= 8'h00;
		14'h167e:	ff_dbi <= 8'h00;
		14'h167f:	ff_dbi <= 8'h00;
		14'h1680:	ff_dbi <= 8'h00;
		14'h1681:	ff_dbi <= 8'h00;
		14'h1682:	ff_dbi <= 8'h00;
		14'h1683:	ff_dbi <= 8'h00;
		14'h1684:	ff_dbi <= 8'h00;
		14'h1685:	ff_dbi <= 8'h00;
		14'h1686:	ff_dbi <= 8'h00;
		14'h1687:	ff_dbi <= 8'h00;
		14'h1688:	ff_dbi <= 8'h00;
		14'h1689:	ff_dbi <= 8'h00;
		14'h168a:	ff_dbi <= 8'h00;
		14'h168b:	ff_dbi <= 8'h00;
		14'h168c:	ff_dbi <= 8'h00;
		14'h168d:	ff_dbi <= 8'h00;
		14'h168e:	ff_dbi <= 8'h00;
		14'h168f:	ff_dbi <= 8'h00;
		14'h1690:	ff_dbi <= 8'h00;
		14'h1691:	ff_dbi <= 8'h00;
		14'h1692:	ff_dbi <= 8'h00;
		14'h1693:	ff_dbi <= 8'h00;
		14'h1694:	ff_dbi <= 8'h00;
		14'h1695:	ff_dbi <= 8'h00;
		14'h1696:	ff_dbi <= 8'h00;
		14'h1697:	ff_dbi <= 8'h00;
		14'h1698:	ff_dbi <= 8'h00;
		14'h1699:	ff_dbi <= 8'h00;
		14'h169a:	ff_dbi <= 8'h00;
		14'h169b:	ff_dbi <= 8'h00;
		14'h169c:	ff_dbi <= 8'h00;
		14'h169d:	ff_dbi <= 8'h00;
		14'h169e:	ff_dbi <= 8'h00;
		14'h169f:	ff_dbi <= 8'h00;
		14'h16a0:	ff_dbi <= 8'h00;
		14'h16a1:	ff_dbi <= 8'h00;
		14'h16a2:	ff_dbi <= 8'h00;
		14'h16a3:	ff_dbi <= 8'h00;
		14'h16a4:	ff_dbi <= 8'h00;
		14'h16a5:	ff_dbi <= 8'h00;
		14'h16a6:	ff_dbi <= 8'h00;
		14'h16a7:	ff_dbi <= 8'h00;
		14'h16a8:	ff_dbi <= 8'h00;
		14'h16a9:	ff_dbi <= 8'h00;
		14'h16aa:	ff_dbi <= 8'h00;
		14'h16ab:	ff_dbi <= 8'h00;
		14'h16ac:	ff_dbi <= 8'h00;
		14'h16ad:	ff_dbi <= 8'h00;
		14'h16ae:	ff_dbi <= 8'h00;
		14'h16af:	ff_dbi <= 8'h00;
		14'h16b0:	ff_dbi <= 8'h00;
		14'h16b1:	ff_dbi <= 8'h00;
		14'h16b2:	ff_dbi <= 8'h00;
		14'h16b3:	ff_dbi <= 8'h00;
		14'h16b4:	ff_dbi <= 8'h00;
		14'h16b5:	ff_dbi <= 8'h00;
		14'h16b6:	ff_dbi <= 8'h00;
		14'h16b7:	ff_dbi <= 8'h00;
		14'h16b8:	ff_dbi <= 8'h00;
		14'h16b9:	ff_dbi <= 8'h00;
		14'h16ba:	ff_dbi <= 8'h00;
		14'h16bb:	ff_dbi <= 8'h00;
		14'h16bc:	ff_dbi <= 8'h00;
		14'h16bd:	ff_dbi <= 8'h00;
		14'h16be:	ff_dbi <= 8'h00;
		14'h16bf:	ff_dbi <= 8'h00;
		14'h16c0:	ff_dbi <= 8'h00;
		14'h16c1:	ff_dbi <= 8'h00;
		14'h16c2:	ff_dbi <= 8'h00;
		14'h16c3:	ff_dbi <= 8'h00;
		14'h16c4:	ff_dbi <= 8'h00;
		14'h16c5:	ff_dbi <= 8'h00;
		14'h16c6:	ff_dbi <= 8'h00;
		14'h16c7:	ff_dbi <= 8'h00;
		14'h16c8:	ff_dbi <= 8'h00;
		14'h16c9:	ff_dbi <= 8'h00;
		14'h16ca:	ff_dbi <= 8'h00;
		14'h16cb:	ff_dbi <= 8'h00;
		14'h16cc:	ff_dbi <= 8'h00;
		14'h16cd:	ff_dbi <= 8'h00;
		14'h16ce:	ff_dbi <= 8'h00;
		14'h16cf:	ff_dbi <= 8'h00;
		14'h16d0:	ff_dbi <= 8'h00;
		14'h16d1:	ff_dbi <= 8'h00;
		14'h16d2:	ff_dbi <= 8'h00;
		14'h16d3:	ff_dbi <= 8'h00;
		14'h16d4:	ff_dbi <= 8'h00;
		14'h16d5:	ff_dbi <= 8'h00;
		14'h16d6:	ff_dbi <= 8'h00;
		14'h16d7:	ff_dbi <= 8'h00;
		14'h16d8:	ff_dbi <= 8'h00;
		14'h16d9:	ff_dbi <= 8'h00;
		14'h16da:	ff_dbi <= 8'h00;
		14'h16db:	ff_dbi <= 8'h00;
		14'h16dc:	ff_dbi <= 8'h00;
		14'h16dd:	ff_dbi <= 8'h00;
		14'h16de:	ff_dbi <= 8'h00;
		14'h16df:	ff_dbi <= 8'h00;
		14'h16e0:	ff_dbi <= 8'h00;
		14'h16e1:	ff_dbi <= 8'h00;
		14'h16e2:	ff_dbi <= 8'h00;
		14'h16e3:	ff_dbi <= 8'h00;
		14'h16e4:	ff_dbi <= 8'h00;
		14'h16e5:	ff_dbi <= 8'h00;
		14'h16e6:	ff_dbi <= 8'h00;
		14'h16e7:	ff_dbi <= 8'h00;
		14'h16e8:	ff_dbi <= 8'h00;
		14'h16e9:	ff_dbi <= 8'h00;
		14'h16ea:	ff_dbi <= 8'h00;
		14'h16eb:	ff_dbi <= 8'h00;
		14'h16ec:	ff_dbi <= 8'h00;
		14'h16ed:	ff_dbi <= 8'h00;
		14'h16ee:	ff_dbi <= 8'h00;
		14'h16ef:	ff_dbi <= 8'h00;
		14'h16f0:	ff_dbi <= 8'h00;
		14'h16f1:	ff_dbi <= 8'h00;
		14'h16f2:	ff_dbi <= 8'h00;
		14'h16f3:	ff_dbi <= 8'h00;
		14'h16f4:	ff_dbi <= 8'h00;
		14'h16f5:	ff_dbi <= 8'h00;
		14'h16f6:	ff_dbi <= 8'h00;
		14'h16f7:	ff_dbi <= 8'h00;
		14'h16f8:	ff_dbi <= 8'h00;
		14'h16f9:	ff_dbi <= 8'h00;
		14'h16fa:	ff_dbi <= 8'h00;
		14'h16fb:	ff_dbi <= 8'h00;
		14'h16fc:	ff_dbi <= 8'h00;
		14'h16fd:	ff_dbi <= 8'h00;
		14'h16fe:	ff_dbi <= 8'h00;
		14'h16ff:	ff_dbi <= 8'h00;
		14'h1700:	ff_dbi <= 8'h00;
		14'h1701:	ff_dbi <= 8'h00;
		14'h1702:	ff_dbi <= 8'h00;
		14'h1703:	ff_dbi <= 8'h00;
		14'h1704:	ff_dbi <= 8'h00;
		14'h1705:	ff_dbi <= 8'h00;
		14'h1706:	ff_dbi <= 8'h00;
		14'h1707:	ff_dbi <= 8'h00;
		14'h1708:	ff_dbi <= 8'h00;
		14'h1709:	ff_dbi <= 8'h00;
		14'h170a:	ff_dbi <= 8'h00;
		14'h170b:	ff_dbi <= 8'h00;
		14'h170c:	ff_dbi <= 8'h00;
		14'h170d:	ff_dbi <= 8'h00;
		14'h170e:	ff_dbi <= 8'h00;
		14'h170f:	ff_dbi <= 8'h00;
		14'h1710:	ff_dbi <= 8'h00;
		14'h1711:	ff_dbi <= 8'h00;
		14'h1712:	ff_dbi <= 8'h00;
		14'h1713:	ff_dbi <= 8'h00;
		14'h1714:	ff_dbi <= 8'h00;
		14'h1715:	ff_dbi <= 8'h00;
		14'h1716:	ff_dbi <= 8'h00;
		14'h1717:	ff_dbi <= 8'h00;
		14'h1718:	ff_dbi <= 8'h00;
		14'h1719:	ff_dbi <= 8'h00;
		14'h171a:	ff_dbi <= 8'h00;
		14'h171b:	ff_dbi <= 8'h00;
		14'h171c:	ff_dbi <= 8'h00;
		14'h171d:	ff_dbi <= 8'h00;
		14'h171e:	ff_dbi <= 8'h00;
		14'h171f:	ff_dbi <= 8'h00;
		14'h1720:	ff_dbi <= 8'h00;
		14'h1721:	ff_dbi <= 8'h00;
		14'h1722:	ff_dbi <= 8'h00;
		14'h1723:	ff_dbi <= 8'h00;
		14'h1724:	ff_dbi <= 8'h00;
		14'h1725:	ff_dbi <= 8'h00;
		14'h1726:	ff_dbi <= 8'h00;
		14'h1727:	ff_dbi <= 8'h00;
		14'h1728:	ff_dbi <= 8'h00;
		14'h1729:	ff_dbi <= 8'h00;
		14'h172a:	ff_dbi <= 8'h00;
		14'h172b:	ff_dbi <= 8'h00;
		14'h172c:	ff_dbi <= 8'h00;
		14'h172d:	ff_dbi <= 8'h00;
		14'h172e:	ff_dbi <= 8'h00;
		14'h172f:	ff_dbi <= 8'h00;
		14'h1730:	ff_dbi <= 8'h00;
		14'h1731:	ff_dbi <= 8'h00;
		14'h1732:	ff_dbi <= 8'h00;
		14'h1733:	ff_dbi <= 8'h00;
		14'h1734:	ff_dbi <= 8'h00;
		14'h1735:	ff_dbi <= 8'h00;
		14'h1736:	ff_dbi <= 8'h00;
		14'h1737:	ff_dbi <= 8'h00;
		14'h1738:	ff_dbi <= 8'h00;
		14'h1739:	ff_dbi <= 8'h00;
		14'h173a:	ff_dbi <= 8'h00;
		14'h173b:	ff_dbi <= 8'h00;
		14'h173c:	ff_dbi <= 8'h00;
		14'h173d:	ff_dbi <= 8'h00;
		14'h173e:	ff_dbi <= 8'h00;
		14'h173f:	ff_dbi <= 8'h00;
		14'h1740:	ff_dbi <= 8'h00;
		14'h1741:	ff_dbi <= 8'h00;
		14'h1742:	ff_dbi <= 8'h00;
		14'h1743:	ff_dbi <= 8'h00;
		14'h1744:	ff_dbi <= 8'h00;
		14'h1745:	ff_dbi <= 8'h00;
		14'h1746:	ff_dbi <= 8'h00;
		14'h1747:	ff_dbi <= 8'h00;
		14'h1748:	ff_dbi <= 8'h00;
		14'h1749:	ff_dbi <= 8'h00;
		14'h174a:	ff_dbi <= 8'h00;
		14'h174b:	ff_dbi <= 8'h00;
		14'h174c:	ff_dbi <= 8'h00;
		14'h174d:	ff_dbi <= 8'h00;
		14'h174e:	ff_dbi <= 8'h00;
		14'h174f:	ff_dbi <= 8'h00;
		14'h1750:	ff_dbi <= 8'h00;
		14'h1751:	ff_dbi <= 8'h00;
		14'h1752:	ff_dbi <= 8'h00;
		14'h1753:	ff_dbi <= 8'h00;
		14'h1754:	ff_dbi <= 8'h00;
		14'h1755:	ff_dbi <= 8'h00;
		14'h1756:	ff_dbi <= 8'h00;
		14'h1757:	ff_dbi <= 8'h00;
		14'h1758:	ff_dbi <= 8'h00;
		14'h1759:	ff_dbi <= 8'h00;
		14'h175a:	ff_dbi <= 8'h00;
		14'h175b:	ff_dbi <= 8'h00;
		14'h175c:	ff_dbi <= 8'h00;
		14'h175d:	ff_dbi <= 8'h00;
		14'h175e:	ff_dbi <= 8'h00;
		14'h175f:	ff_dbi <= 8'h00;
		14'h1760:	ff_dbi <= 8'h00;
		14'h1761:	ff_dbi <= 8'h00;
		14'h1762:	ff_dbi <= 8'h00;
		14'h1763:	ff_dbi <= 8'h00;
		14'h1764:	ff_dbi <= 8'h00;
		14'h1765:	ff_dbi <= 8'h00;
		14'h1766:	ff_dbi <= 8'h00;
		14'h1767:	ff_dbi <= 8'h00;
		14'h1768:	ff_dbi <= 8'h00;
		14'h1769:	ff_dbi <= 8'h00;
		14'h176a:	ff_dbi <= 8'h00;
		14'h176b:	ff_dbi <= 8'h00;
		14'h176c:	ff_dbi <= 8'h00;
		14'h176d:	ff_dbi <= 8'h00;
		14'h176e:	ff_dbi <= 8'h00;
		14'h176f:	ff_dbi <= 8'h00;
		14'h1770:	ff_dbi <= 8'h00;
		14'h1771:	ff_dbi <= 8'h00;
		14'h1772:	ff_dbi <= 8'h00;
		14'h1773:	ff_dbi <= 8'h00;
		14'h1774:	ff_dbi <= 8'h00;
		14'h1775:	ff_dbi <= 8'h00;
		14'h1776:	ff_dbi <= 8'h00;
		14'h1777:	ff_dbi <= 8'h00;
		14'h1778:	ff_dbi <= 8'h00;
		14'h1779:	ff_dbi <= 8'h00;
		14'h177a:	ff_dbi <= 8'h00;
		14'h177b:	ff_dbi <= 8'h00;
		14'h177c:	ff_dbi <= 8'h00;
		14'h177d:	ff_dbi <= 8'h00;
		14'h177e:	ff_dbi <= 8'h00;
		14'h177f:	ff_dbi <= 8'h00;
		14'h1780:	ff_dbi <= 8'h00;
		14'h1781:	ff_dbi <= 8'h00;
		14'h1782:	ff_dbi <= 8'h00;
		14'h1783:	ff_dbi <= 8'h00;
		14'h1784:	ff_dbi <= 8'h00;
		14'h1785:	ff_dbi <= 8'h00;
		14'h1786:	ff_dbi <= 8'h00;
		14'h1787:	ff_dbi <= 8'h00;
		14'h1788:	ff_dbi <= 8'h00;
		14'h1789:	ff_dbi <= 8'h00;
		14'h178a:	ff_dbi <= 8'h00;
		14'h178b:	ff_dbi <= 8'h00;
		14'h178c:	ff_dbi <= 8'h00;
		14'h178d:	ff_dbi <= 8'h00;
		14'h178e:	ff_dbi <= 8'h00;
		14'h178f:	ff_dbi <= 8'h00;
		14'h1790:	ff_dbi <= 8'h00;
		14'h1791:	ff_dbi <= 8'h00;
		14'h1792:	ff_dbi <= 8'h00;
		14'h1793:	ff_dbi <= 8'h00;
		14'h1794:	ff_dbi <= 8'h00;
		14'h1795:	ff_dbi <= 8'h00;
		14'h1796:	ff_dbi <= 8'h00;
		14'h1797:	ff_dbi <= 8'h00;
		14'h1798:	ff_dbi <= 8'h00;
		14'h1799:	ff_dbi <= 8'h00;
		14'h179a:	ff_dbi <= 8'h00;
		14'h179b:	ff_dbi <= 8'h00;
		14'h179c:	ff_dbi <= 8'h00;
		14'h179d:	ff_dbi <= 8'h00;
		14'h179e:	ff_dbi <= 8'h00;
		14'h179f:	ff_dbi <= 8'h00;
		14'h17a0:	ff_dbi <= 8'h00;
		14'h17a1:	ff_dbi <= 8'h00;
		14'h17a2:	ff_dbi <= 8'h00;
		14'h17a3:	ff_dbi <= 8'h00;
		14'h17a4:	ff_dbi <= 8'h00;
		14'h17a5:	ff_dbi <= 8'h00;
		14'h17a6:	ff_dbi <= 8'h00;
		14'h17a7:	ff_dbi <= 8'h00;
		14'h17a8:	ff_dbi <= 8'h00;
		14'h17a9:	ff_dbi <= 8'h00;
		14'h17aa:	ff_dbi <= 8'h00;
		14'h17ab:	ff_dbi <= 8'h00;
		14'h17ac:	ff_dbi <= 8'h00;
		14'h17ad:	ff_dbi <= 8'h00;
		14'h17ae:	ff_dbi <= 8'h00;
		14'h17af:	ff_dbi <= 8'h00;
		14'h17b0:	ff_dbi <= 8'h00;
		14'h17b1:	ff_dbi <= 8'h00;
		14'h17b2:	ff_dbi <= 8'h00;
		14'h17b3:	ff_dbi <= 8'h00;
		14'h17b4:	ff_dbi <= 8'h00;
		14'h17b5:	ff_dbi <= 8'h00;
		14'h17b6:	ff_dbi <= 8'h00;
		14'h17b7:	ff_dbi <= 8'h00;
		14'h17b8:	ff_dbi <= 8'h00;
		14'h17b9:	ff_dbi <= 8'h00;
		14'h17ba:	ff_dbi <= 8'h00;
		14'h17bb:	ff_dbi <= 8'h00;
		14'h17bc:	ff_dbi <= 8'h00;
		14'h17bd:	ff_dbi <= 8'h00;
		14'h17be:	ff_dbi <= 8'h00;
		14'h17bf:	ff_dbi <= 8'h00;
		14'h17c0:	ff_dbi <= 8'h00;
		14'h17c1:	ff_dbi <= 8'h00;
		14'h17c2:	ff_dbi <= 8'h00;
		14'h17c3:	ff_dbi <= 8'h00;
		14'h17c4:	ff_dbi <= 8'h00;
		14'h17c5:	ff_dbi <= 8'h00;
		14'h17c6:	ff_dbi <= 8'h00;
		14'h17c7:	ff_dbi <= 8'h00;
		14'h17c8:	ff_dbi <= 8'h00;
		14'h17c9:	ff_dbi <= 8'h00;
		14'h17ca:	ff_dbi <= 8'h00;
		14'h17cb:	ff_dbi <= 8'h00;
		14'h17cc:	ff_dbi <= 8'h00;
		14'h17cd:	ff_dbi <= 8'h00;
		14'h17ce:	ff_dbi <= 8'h00;
		14'h17cf:	ff_dbi <= 8'h00;
		14'h17d0:	ff_dbi <= 8'h00;
		14'h17d1:	ff_dbi <= 8'h00;
		14'h17d2:	ff_dbi <= 8'h00;
		14'h17d3:	ff_dbi <= 8'h00;
		14'h17d4:	ff_dbi <= 8'h00;
		14'h17d5:	ff_dbi <= 8'h00;
		14'h17d6:	ff_dbi <= 8'h00;
		14'h17d7:	ff_dbi <= 8'h00;
		14'h17d8:	ff_dbi <= 8'h00;
		14'h17d9:	ff_dbi <= 8'h00;
		14'h17da:	ff_dbi <= 8'h00;
		14'h17db:	ff_dbi <= 8'h00;
		14'h17dc:	ff_dbi <= 8'h00;
		14'h17dd:	ff_dbi <= 8'h00;
		14'h17de:	ff_dbi <= 8'h00;
		14'h17df:	ff_dbi <= 8'h00;
		14'h17e0:	ff_dbi <= 8'h00;
		14'h17e1:	ff_dbi <= 8'h00;
		14'h17e2:	ff_dbi <= 8'h00;
		14'h17e3:	ff_dbi <= 8'h00;
		14'h17e4:	ff_dbi <= 8'h00;
		14'h17e5:	ff_dbi <= 8'h00;
		14'h17e6:	ff_dbi <= 8'h00;
		14'h17e7:	ff_dbi <= 8'h00;
		14'h17e8:	ff_dbi <= 8'h00;
		14'h17e9:	ff_dbi <= 8'h00;
		14'h17ea:	ff_dbi <= 8'h00;
		14'h17eb:	ff_dbi <= 8'h00;
		14'h17ec:	ff_dbi <= 8'h00;
		14'h17ed:	ff_dbi <= 8'h00;
		14'h17ee:	ff_dbi <= 8'h00;
		14'h17ef:	ff_dbi <= 8'h00;
		14'h17f0:	ff_dbi <= 8'h00;
		14'h17f1:	ff_dbi <= 8'h00;
		14'h17f2:	ff_dbi <= 8'h00;
		14'h17f3:	ff_dbi <= 8'h00;
		14'h17f4:	ff_dbi <= 8'h00;
		14'h17f5:	ff_dbi <= 8'h00;
		14'h17f6:	ff_dbi <= 8'h00;
		14'h17f7:	ff_dbi <= 8'h00;
		14'h17f8:	ff_dbi <= 8'h00;
		14'h17f9:	ff_dbi <= 8'h00;
		14'h17fa:	ff_dbi <= 8'h00;
		14'h17fb:	ff_dbi <= 8'h00;
		14'h17fc:	ff_dbi <= 8'h00;
		14'h17fd:	ff_dbi <= 8'h00;
		14'h17fe:	ff_dbi <= 8'h00;
		14'h17ff:	ff_dbi <= 8'h00;
		14'h1800:	ff_dbi <= 8'h20;
		14'h1801:	ff_dbi <= 8'h20;
		14'h1802:	ff_dbi <= 8'h4d;
		14'h1803:	ff_dbi <= 8'h53;
		14'h1804:	ff_dbi <= 8'h58;
		14'h1805:	ff_dbi <= 8'h20;
		14'h1806:	ff_dbi <= 8'h42;
		14'h1807:	ff_dbi <= 8'h41;
		14'h1808:	ff_dbi <= 8'h53;
		14'h1809:	ff_dbi <= 8'h49;
		14'h180a:	ff_dbi <= 8'h43;
		14'h180b:	ff_dbi <= 8'h20;
		14'h180c:	ff_dbi <= 8'h76;
		14'h180d:	ff_dbi <= 8'h65;
		14'h180e:	ff_dbi <= 8'h72;
		14'h180f:	ff_dbi <= 8'h73;
		14'h1810:	ff_dbi <= 8'h69;
		14'h1811:	ff_dbi <= 8'h6f;
		14'h1812:	ff_dbi <= 8'h6e;
		14'h1813:	ff_dbi <= 8'h20;
		14'h1814:	ff_dbi <= 8'h34;
		14'h1815:	ff_dbi <= 8'h2e;
		14'h1816:	ff_dbi <= 8'h31;
		14'h1817:	ff_dbi <= 8'h20;
		14'h1818:	ff_dbi <= 8'h20;
		14'h1819:	ff_dbi <= 8'h20;
		14'h181a:	ff_dbi <= 8'h20;
		14'h181b:	ff_dbi <= 8'h20;
		14'h181c:	ff_dbi <= 8'h20;
		14'h181d:	ff_dbi <= 8'h20;
		14'h181e:	ff_dbi <= 8'h20;
		14'h181f:	ff_dbi <= 8'h20;
		14'h1820:	ff_dbi <= 8'h20;
		14'h1821:	ff_dbi <= 8'h20;
		14'h1822:	ff_dbi <= 8'h43;
		14'h1823:	ff_dbi <= 8'h6f;
		14'h1824:	ff_dbi <= 8'h70;
		14'h1825:	ff_dbi <= 8'h79;
		14'h1826:	ff_dbi <= 8'h72;
		14'h1827:	ff_dbi <= 8'h69;
		14'h1828:	ff_dbi <= 8'h67;
		14'h1829:	ff_dbi <= 8'h68;
		14'h182a:	ff_dbi <= 8'h74;
		14'h182b:	ff_dbi <= 8'h20;
		14'h182c:	ff_dbi <= 8'h31;
		14'h182d:	ff_dbi <= 8'h39;
		14'h182e:	ff_dbi <= 8'h39;
		14'h182f:	ff_dbi <= 8'h30;
		14'h1830:	ff_dbi <= 8'h20;
		14'h1831:	ff_dbi <= 8'h62;
		14'h1832:	ff_dbi <= 8'h79;
		14'h1833:	ff_dbi <= 8'h20;
		14'h1834:	ff_dbi <= 8'h4d;
		14'h1835:	ff_dbi <= 8'h69;
		14'h1836:	ff_dbi <= 8'h63;
		14'h1837:	ff_dbi <= 8'h72;
		14'h1838:	ff_dbi <= 8'h6f;
		14'h1839:	ff_dbi <= 8'h73;
		14'h183a:	ff_dbi <= 8'h6f;
		14'h183b:	ff_dbi <= 8'h66;
		14'h183c:	ff_dbi <= 8'h74;
		14'h183d:	ff_dbi <= 8'h20;
		14'h183e:	ff_dbi <= 8'h20;
		14'h183f:	ff_dbi <= 8'h20;
		14'h1840:	ff_dbi <= 8'h20;
		14'h1841:	ff_dbi <= 8'h20;
		14'h1842:	ff_dbi <= 8'h32;
		14'h1843:	ff_dbi <= 8'h35;
		14'h1844:	ff_dbi <= 8'h32;
		14'h1845:	ff_dbi <= 8'h37;
		14'h1846:	ff_dbi <= 8'h31;
		14'h1847:	ff_dbi <= 8'h20;
		14'h1848:	ff_dbi <= 8'h42;
		14'h1849:	ff_dbi <= 8'h79;
		14'h184a:	ff_dbi <= 8'h74;
		14'h184b:	ff_dbi <= 8'h65;
		14'h184c:	ff_dbi <= 8'h73;
		14'h184d:	ff_dbi <= 8'h20;
		14'h184e:	ff_dbi <= 8'h66;
		14'h184f:	ff_dbi <= 8'h72;
		14'h1850:	ff_dbi <= 8'h65;
		14'h1851:	ff_dbi <= 8'h65;
		14'h1852:	ff_dbi <= 8'h20;
		14'h1853:	ff_dbi <= 8'h20;
		14'h1854:	ff_dbi <= 8'h20;
		14'h1855:	ff_dbi <= 8'h20;
		14'h1856:	ff_dbi <= 8'h20;
		14'h1857:	ff_dbi <= 8'h20;
		14'h1858:	ff_dbi <= 8'h20;
		14'h1859:	ff_dbi <= 8'h20;
		14'h185a:	ff_dbi <= 8'h20;
		14'h185b:	ff_dbi <= 8'h20;
		14'h185c:	ff_dbi <= 8'h20;
		14'h185d:	ff_dbi <= 8'h20;
		14'h185e:	ff_dbi <= 8'h20;
		14'h185f:	ff_dbi <= 8'h20;
		14'h1860:	ff_dbi <= 8'h20;
		14'h1861:	ff_dbi <= 8'h20;
		14'h1862:	ff_dbi <= 8'h44;
		14'h1863:	ff_dbi <= 8'h69;
		14'h1864:	ff_dbi <= 8'h73;
		14'h1865:	ff_dbi <= 8'h6b;
		14'h1866:	ff_dbi <= 8'h20;
		14'h1867:	ff_dbi <= 8'h42;
		14'h1868:	ff_dbi <= 8'h41;
		14'h1869:	ff_dbi <= 8'h53;
		14'h186a:	ff_dbi <= 8'h49;
		14'h186b:	ff_dbi <= 8'h43;
		14'h186c:	ff_dbi <= 8'h20;
		14'h186d:	ff_dbi <= 8'h76;
		14'h186e:	ff_dbi <= 8'h65;
		14'h186f:	ff_dbi <= 8'h72;
		14'h1870:	ff_dbi <= 8'h73;
		14'h1871:	ff_dbi <= 8'h69;
		14'h1872:	ff_dbi <= 8'h6f;
		14'h1873:	ff_dbi <= 8'h6e;
		14'h1874:	ff_dbi <= 8'h20;
		14'h1875:	ff_dbi <= 8'h32;
		14'h1876:	ff_dbi <= 8'h2e;
		14'h1877:	ff_dbi <= 8'h30;
		14'h1878:	ff_dbi <= 8'h31;
		14'h1879:	ff_dbi <= 8'h20;
		14'h187a:	ff_dbi <= 8'h20;
		14'h187b:	ff_dbi <= 8'h20;
		14'h187c:	ff_dbi <= 8'h20;
		14'h187d:	ff_dbi <= 8'h20;
		14'h187e:	ff_dbi <= 8'h20;
		14'h187f:	ff_dbi <= 8'h20;
		14'h1880:	ff_dbi <= 8'h20;
		14'h1881:	ff_dbi <= 8'h20;
		14'h1882:	ff_dbi <= 8'h4f;
		14'h1883:	ff_dbi <= 8'h6b;
		14'h1884:	ff_dbi <= 8'h20;
		14'h1885:	ff_dbi <= 8'h20;
		14'h1886:	ff_dbi <= 8'h20;
		14'h1887:	ff_dbi <= 8'h20;
		14'h1888:	ff_dbi <= 8'h20;
		14'h1889:	ff_dbi <= 8'h20;
		14'h188a:	ff_dbi <= 8'h20;
		14'h188b:	ff_dbi <= 8'h20;
		14'h188c:	ff_dbi <= 8'h20;
		14'h188d:	ff_dbi <= 8'h20;
		14'h188e:	ff_dbi <= 8'h20;
		14'h188f:	ff_dbi <= 8'h20;
		14'h1890:	ff_dbi <= 8'h20;
		14'h1891:	ff_dbi <= 8'h20;
		14'h1892:	ff_dbi <= 8'h20;
		14'h1893:	ff_dbi <= 8'h20;
		14'h1894:	ff_dbi <= 8'h20;
		14'h1895:	ff_dbi <= 8'h20;
		14'h1896:	ff_dbi <= 8'h20;
		14'h1897:	ff_dbi <= 8'h20;
		14'h1898:	ff_dbi <= 8'h20;
		14'h1899:	ff_dbi <= 8'h20;
		14'h189a:	ff_dbi <= 8'h20;
		14'h189b:	ff_dbi <= 8'h20;
		14'h189c:	ff_dbi <= 8'h20;
		14'h189d:	ff_dbi <= 8'h20;
		14'h189e:	ff_dbi <= 8'h20;
		14'h189f:	ff_dbi <= 8'h20;
		14'h18a0:	ff_dbi <= 8'h20;
		14'h18a1:	ff_dbi <= 8'h20;
		14'h18a2:	ff_dbi <= 8'hff;
		14'h18a3:	ff_dbi <= 8'h20;
		14'h18a4:	ff_dbi <= 8'h20;
		14'h18a5:	ff_dbi <= 8'h20;
		14'h18a6:	ff_dbi <= 8'h20;
		14'h18a7:	ff_dbi <= 8'h20;
		14'h18a8:	ff_dbi <= 8'h20;
		14'h18a9:	ff_dbi <= 8'h20;
		14'h18aa:	ff_dbi <= 8'h20;
		14'h18ab:	ff_dbi <= 8'h20;
		14'h18ac:	ff_dbi <= 8'h20;
		14'h18ad:	ff_dbi <= 8'h20;
		14'h18ae:	ff_dbi <= 8'h20;
		14'h18af:	ff_dbi <= 8'h20;
		14'h18b0:	ff_dbi <= 8'h20;
		14'h18b1:	ff_dbi <= 8'h20;
		14'h18b2:	ff_dbi <= 8'h20;
		14'h18b3:	ff_dbi <= 8'h20;
		14'h18b4:	ff_dbi <= 8'h20;
		14'h18b5:	ff_dbi <= 8'h20;
		14'h18b6:	ff_dbi <= 8'h20;
		14'h18b7:	ff_dbi <= 8'h20;
		14'h18b8:	ff_dbi <= 8'h20;
		14'h18b9:	ff_dbi <= 8'h20;
		14'h18ba:	ff_dbi <= 8'h20;
		14'h18bb:	ff_dbi <= 8'h20;
		14'h18bc:	ff_dbi <= 8'h20;
		14'h18bd:	ff_dbi <= 8'h20;
		14'h18be:	ff_dbi <= 8'h20;
		14'h18bf:	ff_dbi <= 8'h20;
		14'h18c0:	ff_dbi <= 8'h20;
		14'h18c1:	ff_dbi <= 8'h20;
		14'h18c2:	ff_dbi <= 8'h20;
		14'h18c3:	ff_dbi <= 8'h20;
		14'h18c4:	ff_dbi <= 8'h20;
		14'h18c5:	ff_dbi <= 8'h20;
		14'h18c6:	ff_dbi <= 8'h20;
		14'h18c7:	ff_dbi <= 8'h20;
		14'h18c8:	ff_dbi <= 8'h20;
		14'h18c9:	ff_dbi <= 8'h20;
		14'h18ca:	ff_dbi <= 8'h20;
		14'h18cb:	ff_dbi <= 8'h20;
		14'h18cc:	ff_dbi <= 8'h20;
		14'h18cd:	ff_dbi <= 8'h20;
		14'h18ce:	ff_dbi <= 8'h20;
		14'h18cf:	ff_dbi <= 8'h20;
		14'h18d0:	ff_dbi <= 8'h20;
		14'h18d1:	ff_dbi <= 8'h20;
		14'h18d2:	ff_dbi <= 8'h20;
		14'h18d3:	ff_dbi <= 8'h20;
		14'h18d4:	ff_dbi <= 8'h20;
		14'h18d5:	ff_dbi <= 8'h20;
		14'h18d6:	ff_dbi <= 8'h20;
		14'h18d7:	ff_dbi <= 8'h20;
		14'h18d8:	ff_dbi <= 8'h20;
		14'h18d9:	ff_dbi <= 8'h20;
		14'h18da:	ff_dbi <= 8'h20;
		14'h18db:	ff_dbi <= 8'h20;
		14'h18dc:	ff_dbi <= 8'h20;
		14'h18dd:	ff_dbi <= 8'h20;
		14'h18de:	ff_dbi <= 8'h20;
		14'h18df:	ff_dbi <= 8'h20;
		14'h18e0:	ff_dbi <= 8'h20;
		14'h18e1:	ff_dbi <= 8'h20;
		14'h18e2:	ff_dbi <= 8'h20;
		14'h18e3:	ff_dbi <= 8'h20;
		14'h18e4:	ff_dbi <= 8'h20;
		14'h18e5:	ff_dbi <= 8'h20;
		14'h18e6:	ff_dbi <= 8'h20;
		14'h18e7:	ff_dbi <= 8'h20;
		14'h18e8:	ff_dbi <= 8'h20;
		14'h18e9:	ff_dbi <= 8'h20;
		14'h18ea:	ff_dbi <= 8'h20;
		14'h18eb:	ff_dbi <= 8'h20;
		14'h18ec:	ff_dbi <= 8'h20;
		14'h18ed:	ff_dbi <= 8'h20;
		14'h18ee:	ff_dbi <= 8'h20;
		14'h18ef:	ff_dbi <= 8'h20;
		14'h18f0:	ff_dbi <= 8'h20;
		14'h18f1:	ff_dbi <= 8'h20;
		14'h18f2:	ff_dbi <= 8'h20;
		14'h18f3:	ff_dbi <= 8'h20;
		14'h18f4:	ff_dbi <= 8'h20;
		14'h18f5:	ff_dbi <= 8'h20;
		14'h18f6:	ff_dbi <= 8'h20;
		14'h18f7:	ff_dbi <= 8'h20;
		14'h18f8:	ff_dbi <= 8'h20;
		14'h18f9:	ff_dbi <= 8'h20;
		14'h18fa:	ff_dbi <= 8'h20;
		14'h18fb:	ff_dbi <= 8'h20;
		14'h18fc:	ff_dbi <= 8'h20;
		14'h18fd:	ff_dbi <= 8'h20;
		14'h18fe:	ff_dbi <= 8'h20;
		14'h18ff:	ff_dbi <= 8'h20;
		14'h1900:	ff_dbi <= 8'h20;
		14'h1901:	ff_dbi <= 8'h20;
		14'h1902:	ff_dbi <= 8'h20;
		14'h1903:	ff_dbi <= 8'h20;
		14'h1904:	ff_dbi <= 8'h20;
		14'h1905:	ff_dbi <= 8'h20;
		14'h1906:	ff_dbi <= 8'h20;
		14'h1907:	ff_dbi <= 8'h20;
		14'h1908:	ff_dbi <= 8'h20;
		14'h1909:	ff_dbi <= 8'h20;
		14'h190a:	ff_dbi <= 8'h20;
		14'h190b:	ff_dbi <= 8'h20;
		14'h190c:	ff_dbi <= 8'h20;
		14'h190d:	ff_dbi <= 8'h20;
		14'h190e:	ff_dbi <= 8'h20;
		14'h190f:	ff_dbi <= 8'h20;
		14'h1910:	ff_dbi <= 8'h20;
		14'h1911:	ff_dbi <= 8'h20;
		14'h1912:	ff_dbi <= 8'h20;
		14'h1913:	ff_dbi <= 8'h20;
		14'h1914:	ff_dbi <= 8'h20;
		14'h1915:	ff_dbi <= 8'h20;
		14'h1916:	ff_dbi <= 8'h20;
		14'h1917:	ff_dbi <= 8'h20;
		14'h1918:	ff_dbi <= 8'h20;
		14'h1919:	ff_dbi <= 8'h20;
		14'h191a:	ff_dbi <= 8'h20;
		14'h191b:	ff_dbi <= 8'h20;
		14'h191c:	ff_dbi <= 8'h20;
		14'h191d:	ff_dbi <= 8'h20;
		14'h191e:	ff_dbi <= 8'h20;
		14'h191f:	ff_dbi <= 8'h20;
		14'h1920:	ff_dbi <= 8'h20;
		14'h1921:	ff_dbi <= 8'h20;
		14'h1922:	ff_dbi <= 8'h20;
		14'h1923:	ff_dbi <= 8'h20;
		14'h1924:	ff_dbi <= 8'h20;
		14'h1925:	ff_dbi <= 8'h20;
		14'h1926:	ff_dbi <= 8'h20;
		14'h1927:	ff_dbi <= 8'h20;
		14'h1928:	ff_dbi <= 8'h20;
		14'h1929:	ff_dbi <= 8'h20;
		14'h192a:	ff_dbi <= 8'h20;
		14'h192b:	ff_dbi <= 8'h20;
		14'h192c:	ff_dbi <= 8'h20;
		14'h192d:	ff_dbi <= 8'h20;
		14'h192e:	ff_dbi <= 8'h20;
		14'h192f:	ff_dbi <= 8'h20;
		14'h1930:	ff_dbi <= 8'h20;
		14'h1931:	ff_dbi <= 8'h20;
		14'h1932:	ff_dbi <= 8'h20;
		14'h1933:	ff_dbi <= 8'h20;
		14'h1934:	ff_dbi <= 8'h20;
		14'h1935:	ff_dbi <= 8'h20;
		14'h1936:	ff_dbi <= 8'h20;
		14'h1937:	ff_dbi <= 8'h20;
		14'h1938:	ff_dbi <= 8'h20;
		14'h1939:	ff_dbi <= 8'h20;
		14'h193a:	ff_dbi <= 8'h20;
		14'h193b:	ff_dbi <= 8'h20;
		14'h193c:	ff_dbi <= 8'h20;
		14'h193d:	ff_dbi <= 8'h20;
		14'h193e:	ff_dbi <= 8'h20;
		14'h193f:	ff_dbi <= 8'h20;
		14'h1940:	ff_dbi <= 8'h20;
		14'h1941:	ff_dbi <= 8'h20;
		14'h1942:	ff_dbi <= 8'h20;
		14'h1943:	ff_dbi <= 8'h20;
		14'h1944:	ff_dbi <= 8'h20;
		14'h1945:	ff_dbi <= 8'h20;
		14'h1946:	ff_dbi <= 8'h20;
		14'h1947:	ff_dbi <= 8'h20;
		14'h1948:	ff_dbi <= 8'h20;
		14'h1949:	ff_dbi <= 8'h20;
		14'h194a:	ff_dbi <= 8'h20;
		14'h194b:	ff_dbi <= 8'h20;
		14'h194c:	ff_dbi <= 8'h20;
		14'h194d:	ff_dbi <= 8'h20;
		14'h194e:	ff_dbi <= 8'h20;
		14'h194f:	ff_dbi <= 8'h20;
		14'h1950:	ff_dbi <= 8'h20;
		14'h1951:	ff_dbi <= 8'h20;
		14'h1952:	ff_dbi <= 8'h20;
		14'h1953:	ff_dbi <= 8'h20;
		14'h1954:	ff_dbi <= 8'h20;
		14'h1955:	ff_dbi <= 8'h20;
		14'h1956:	ff_dbi <= 8'h20;
		14'h1957:	ff_dbi <= 8'h20;
		14'h1958:	ff_dbi <= 8'h20;
		14'h1959:	ff_dbi <= 8'h20;
		14'h195a:	ff_dbi <= 8'h20;
		14'h195b:	ff_dbi <= 8'h20;
		14'h195c:	ff_dbi <= 8'h20;
		14'h195d:	ff_dbi <= 8'h20;
		14'h195e:	ff_dbi <= 8'h20;
		14'h195f:	ff_dbi <= 8'h20;
		14'h1960:	ff_dbi <= 8'h20;
		14'h1961:	ff_dbi <= 8'h20;
		14'h1962:	ff_dbi <= 8'h20;
		14'h1963:	ff_dbi <= 8'h20;
		14'h1964:	ff_dbi <= 8'h20;
		14'h1965:	ff_dbi <= 8'h20;
		14'h1966:	ff_dbi <= 8'h20;
		14'h1967:	ff_dbi <= 8'h20;
		14'h1968:	ff_dbi <= 8'h20;
		14'h1969:	ff_dbi <= 8'h20;
		14'h196a:	ff_dbi <= 8'h20;
		14'h196b:	ff_dbi <= 8'h20;
		14'h196c:	ff_dbi <= 8'h20;
		14'h196d:	ff_dbi <= 8'h20;
		14'h196e:	ff_dbi <= 8'h20;
		14'h196f:	ff_dbi <= 8'h20;
		14'h1970:	ff_dbi <= 8'h20;
		14'h1971:	ff_dbi <= 8'h20;
		14'h1972:	ff_dbi <= 8'h20;
		14'h1973:	ff_dbi <= 8'h20;
		14'h1974:	ff_dbi <= 8'h20;
		14'h1975:	ff_dbi <= 8'h20;
		14'h1976:	ff_dbi <= 8'h20;
		14'h1977:	ff_dbi <= 8'h20;
		14'h1978:	ff_dbi <= 8'h20;
		14'h1979:	ff_dbi <= 8'h20;
		14'h197a:	ff_dbi <= 8'h20;
		14'h197b:	ff_dbi <= 8'h20;
		14'h197c:	ff_dbi <= 8'h20;
		14'h197d:	ff_dbi <= 8'h20;
		14'h197e:	ff_dbi <= 8'h20;
		14'h197f:	ff_dbi <= 8'h20;
		14'h1980:	ff_dbi <= 8'h20;
		14'h1981:	ff_dbi <= 8'h20;
		14'h1982:	ff_dbi <= 8'h20;
		14'h1983:	ff_dbi <= 8'h20;
		14'h1984:	ff_dbi <= 8'h20;
		14'h1985:	ff_dbi <= 8'h20;
		14'h1986:	ff_dbi <= 8'h20;
		14'h1987:	ff_dbi <= 8'h20;
		14'h1988:	ff_dbi <= 8'h20;
		14'h1989:	ff_dbi <= 8'h20;
		14'h198a:	ff_dbi <= 8'h20;
		14'h198b:	ff_dbi <= 8'h20;
		14'h198c:	ff_dbi <= 8'h20;
		14'h198d:	ff_dbi <= 8'h20;
		14'h198e:	ff_dbi <= 8'h20;
		14'h198f:	ff_dbi <= 8'h20;
		14'h1990:	ff_dbi <= 8'h20;
		14'h1991:	ff_dbi <= 8'h20;
		14'h1992:	ff_dbi <= 8'h20;
		14'h1993:	ff_dbi <= 8'h20;
		14'h1994:	ff_dbi <= 8'h20;
		14'h1995:	ff_dbi <= 8'h20;
		14'h1996:	ff_dbi <= 8'h20;
		14'h1997:	ff_dbi <= 8'h20;
		14'h1998:	ff_dbi <= 8'h20;
		14'h1999:	ff_dbi <= 8'h20;
		14'h199a:	ff_dbi <= 8'h20;
		14'h199b:	ff_dbi <= 8'h20;
		14'h199c:	ff_dbi <= 8'h20;
		14'h199d:	ff_dbi <= 8'h20;
		14'h199e:	ff_dbi <= 8'h20;
		14'h199f:	ff_dbi <= 8'h20;
		14'h19a0:	ff_dbi <= 8'h20;
		14'h19a1:	ff_dbi <= 8'h20;
		14'h19a2:	ff_dbi <= 8'h20;
		14'h19a3:	ff_dbi <= 8'h20;
		14'h19a4:	ff_dbi <= 8'h20;
		14'h19a5:	ff_dbi <= 8'h20;
		14'h19a6:	ff_dbi <= 8'h20;
		14'h19a7:	ff_dbi <= 8'h20;
		14'h19a8:	ff_dbi <= 8'h20;
		14'h19a9:	ff_dbi <= 8'h20;
		14'h19aa:	ff_dbi <= 8'h20;
		14'h19ab:	ff_dbi <= 8'h20;
		14'h19ac:	ff_dbi <= 8'h20;
		14'h19ad:	ff_dbi <= 8'h20;
		14'h19ae:	ff_dbi <= 8'h20;
		14'h19af:	ff_dbi <= 8'h20;
		14'h19b0:	ff_dbi <= 8'h20;
		14'h19b1:	ff_dbi <= 8'h20;
		14'h19b2:	ff_dbi <= 8'h20;
		14'h19b3:	ff_dbi <= 8'h20;
		14'h19b4:	ff_dbi <= 8'h20;
		14'h19b5:	ff_dbi <= 8'h20;
		14'h19b6:	ff_dbi <= 8'h20;
		14'h19b7:	ff_dbi <= 8'h20;
		14'h19b8:	ff_dbi <= 8'h20;
		14'h19b9:	ff_dbi <= 8'h20;
		14'h19ba:	ff_dbi <= 8'h20;
		14'h19bb:	ff_dbi <= 8'h20;
		14'h19bc:	ff_dbi <= 8'h20;
		14'h19bd:	ff_dbi <= 8'h20;
		14'h19be:	ff_dbi <= 8'h20;
		14'h19bf:	ff_dbi <= 8'h20;
		14'h19c0:	ff_dbi <= 8'h20;
		14'h19c1:	ff_dbi <= 8'h20;
		14'h19c2:	ff_dbi <= 8'h20;
		14'h19c3:	ff_dbi <= 8'h20;
		14'h19c4:	ff_dbi <= 8'h20;
		14'h19c5:	ff_dbi <= 8'h20;
		14'h19c6:	ff_dbi <= 8'h20;
		14'h19c7:	ff_dbi <= 8'h20;
		14'h19c8:	ff_dbi <= 8'h20;
		14'h19c9:	ff_dbi <= 8'h20;
		14'h19ca:	ff_dbi <= 8'h20;
		14'h19cb:	ff_dbi <= 8'h20;
		14'h19cc:	ff_dbi <= 8'h20;
		14'h19cd:	ff_dbi <= 8'h20;
		14'h19ce:	ff_dbi <= 8'h20;
		14'h19cf:	ff_dbi <= 8'h20;
		14'h19d0:	ff_dbi <= 8'h20;
		14'h19d1:	ff_dbi <= 8'h20;
		14'h19d2:	ff_dbi <= 8'h20;
		14'h19d3:	ff_dbi <= 8'h20;
		14'h19d4:	ff_dbi <= 8'h20;
		14'h19d5:	ff_dbi <= 8'h20;
		14'h19d6:	ff_dbi <= 8'h20;
		14'h19d7:	ff_dbi <= 8'h20;
		14'h19d8:	ff_dbi <= 8'h20;
		14'h19d9:	ff_dbi <= 8'h20;
		14'h19da:	ff_dbi <= 8'h20;
		14'h19db:	ff_dbi <= 8'h20;
		14'h19dc:	ff_dbi <= 8'h20;
		14'h19dd:	ff_dbi <= 8'h20;
		14'h19de:	ff_dbi <= 8'h20;
		14'h19df:	ff_dbi <= 8'h20;
		14'h19e0:	ff_dbi <= 8'h20;
		14'h19e1:	ff_dbi <= 8'h20;
		14'h19e2:	ff_dbi <= 8'h20;
		14'h19e3:	ff_dbi <= 8'h20;
		14'h19e4:	ff_dbi <= 8'h20;
		14'h19e5:	ff_dbi <= 8'h20;
		14'h19e6:	ff_dbi <= 8'h20;
		14'h19e7:	ff_dbi <= 8'h20;
		14'h19e8:	ff_dbi <= 8'h20;
		14'h19e9:	ff_dbi <= 8'h20;
		14'h19ea:	ff_dbi <= 8'h20;
		14'h19eb:	ff_dbi <= 8'h20;
		14'h19ec:	ff_dbi <= 8'h20;
		14'h19ed:	ff_dbi <= 8'h20;
		14'h19ee:	ff_dbi <= 8'h20;
		14'h19ef:	ff_dbi <= 8'h20;
		14'h19f0:	ff_dbi <= 8'h20;
		14'h19f1:	ff_dbi <= 8'h20;
		14'h19f2:	ff_dbi <= 8'h20;
		14'h19f3:	ff_dbi <= 8'h20;
		14'h19f4:	ff_dbi <= 8'h20;
		14'h19f5:	ff_dbi <= 8'h20;
		14'h19f6:	ff_dbi <= 8'h20;
		14'h19f7:	ff_dbi <= 8'h20;
		14'h19f8:	ff_dbi <= 8'h20;
		14'h19f9:	ff_dbi <= 8'h20;
		14'h19fa:	ff_dbi <= 8'h20;
		14'h19fb:	ff_dbi <= 8'h20;
		14'h19fc:	ff_dbi <= 8'h20;
		14'h19fd:	ff_dbi <= 8'h20;
		14'h19fe:	ff_dbi <= 8'h20;
		14'h19ff:	ff_dbi <= 8'h20;
		14'h1a00:	ff_dbi <= 8'h20;
		14'h1a01:	ff_dbi <= 8'h20;
		14'h1a02:	ff_dbi <= 8'h20;
		14'h1a03:	ff_dbi <= 8'h20;
		14'h1a04:	ff_dbi <= 8'h20;
		14'h1a05:	ff_dbi <= 8'h20;
		14'h1a06:	ff_dbi <= 8'h20;
		14'h1a07:	ff_dbi <= 8'h20;
		14'h1a08:	ff_dbi <= 8'h20;
		14'h1a09:	ff_dbi <= 8'h20;
		14'h1a0a:	ff_dbi <= 8'h20;
		14'h1a0b:	ff_dbi <= 8'h20;
		14'h1a0c:	ff_dbi <= 8'h20;
		14'h1a0d:	ff_dbi <= 8'h20;
		14'h1a0e:	ff_dbi <= 8'h20;
		14'h1a0f:	ff_dbi <= 8'h20;
		14'h1a10:	ff_dbi <= 8'h20;
		14'h1a11:	ff_dbi <= 8'h20;
		14'h1a12:	ff_dbi <= 8'h20;
		14'h1a13:	ff_dbi <= 8'h20;
		14'h1a14:	ff_dbi <= 8'h20;
		14'h1a15:	ff_dbi <= 8'h20;
		14'h1a16:	ff_dbi <= 8'h20;
		14'h1a17:	ff_dbi <= 8'h20;
		14'h1a18:	ff_dbi <= 8'h20;
		14'h1a19:	ff_dbi <= 8'h20;
		14'h1a1a:	ff_dbi <= 8'h20;
		14'h1a1b:	ff_dbi <= 8'h20;
		14'h1a1c:	ff_dbi <= 8'h20;
		14'h1a1d:	ff_dbi <= 8'h20;
		14'h1a1e:	ff_dbi <= 8'h20;
		14'h1a1f:	ff_dbi <= 8'h20;
		14'h1a20:	ff_dbi <= 8'h20;
		14'h1a21:	ff_dbi <= 8'h20;
		14'h1a22:	ff_dbi <= 8'h20;
		14'h1a23:	ff_dbi <= 8'h20;
		14'h1a24:	ff_dbi <= 8'h20;
		14'h1a25:	ff_dbi <= 8'h20;
		14'h1a26:	ff_dbi <= 8'h20;
		14'h1a27:	ff_dbi <= 8'h20;
		14'h1a28:	ff_dbi <= 8'h20;
		14'h1a29:	ff_dbi <= 8'h20;
		14'h1a2a:	ff_dbi <= 8'h20;
		14'h1a2b:	ff_dbi <= 8'h20;
		14'h1a2c:	ff_dbi <= 8'h20;
		14'h1a2d:	ff_dbi <= 8'h20;
		14'h1a2e:	ff_dbi <= 8'h20;
		14'h1a2f:	ff_dbi <= 8'h20;
		14'h1a30:	ff_dbi <= 8'h20;
		14'h1a31:	ff_dbi <= 8'h20;
		14'h1a32:	ff_dbi <= 8'h20;
		14'h1a33:	ff_dbi <= 8'h20;
		14'h1a34:	ff_dbi <= 8'h20;
		14'h1a35:	ff_dbi <= 8'h20;
		14'h1a36:	ff_dbi <= 8'h20;
		14'h1a37:	ff_dbi <= 8'h20;
		14'h1a38:	ff_dbi <= 8'h20;
		14'h1a39:	ff_dbi <= 8'h20;
		14'h1a3a:	ff_dbi <= 8'h20;
		14'h1a3b:	ff_dbi <= 8'h20;
		14'h1a3c:	ff_dbi <= 8'h20;
		14'h1a3d:	ff_dbi <= 8'h20;
		14'h1a3e:	ff_dbi <= 8'h20;
		14'h1a3f:	ff_dbi <= 8'h20;
		14'h1a40:	ff_dbi <= 8'h20;
		14'h1a41:	ff_dbi <= 8'h20;
		14'h1a42:	ff_dbi <= 8'h20;
		14'h1a43:	ff_dbi <= 8'h20;
		14'h1a44:	ff_dbi <= 8'h20;
		14'h1a45:	ff_dbi <= 8'h20;
		14'h1a46:	ff_dbi <= 8'h20;
		14'h1a47:	ff_dbi <= 8'h20;
		14'h1a48:	ff_dbi <= 8'h20;
		14'h1a49:	ff_dbi <= 8'h20;
		14'h1a4a:	ff_dbi <= 8'h20;
		14'h1a4b:	ff_dbi <= 8'h20;
		14'h1a4c:	ff_dbi <= 8'h20;
		14'h1a4d:	ff_dbi <= 8'h20;
		14'h1a4e:	ff_dbi <= 8'h20;
		14'h1a4f:	ff_dbi <= 8'h20;
		14'h1a50:	ff_dbi <= 8'h20;
		14'h1a51:	ff_dbi <= 8'h20;
		14'h1a52:	ff_dbi <= 8'h20;
		14'h1a53:	ff_dbi <= 8'h20;
		14'h1a54:	ff_dbi <= 8'h20;
		14'h1a55:	ff_dbi <= 8'h20;
		14'h1a56:	ff_dbi <= 8'h20;
		14'h1a57:	ff_dbi <= 8'h20;
		14'h1a58:	ff_dbi <= 8'h20;
		14'h1a59:	ff_dbi <= 8'h20;
		14'h1a5a:	ff_dbi <= 8'h20;
		14'h1a5b:	ff_dbi <= 8'h20;
		14'h1a5c:	ff_dbi <= 8'h20;
		14'h1a5d:	ff_dbi <= 8'h20;
		14'h1a5e:	ff_dbi <= 8'h20;
		14'h1a5f:	ff_dbi <= 8'h20;
		14'h1a60:	ff_dbi <= 8'h20;
		14'h1a61:	ff_dbi <= 8'h20;
		14'h1a62:	ff_dbi <= 8'h20;
		14'h1a63:	ff_dbi <= 8'h20;
		14'h1a64:	ff_dbi <= 8'h20;
		14'h1a65:	ff_dbi <= 8'h20;
		14'h1a66:	ff_dbi <= 8'h20;
		14'h1a67:	ff_dbi <= 8'h20;
		14'h1a68:	ff_dbi <= 8'h20;
		14'h1a69:	ff_dbi <= 8'h20;
		14'h1a6a:	ff_dbi <= 8'h20;
		14'h1a6b:	ff_dbi <= 8'h20;
		14'h1a6c:	ff_dbi <= 8'h20;
		14'h1a6d:	ff_dbi <= 8'h20;
		14'h1a6e:	ff_dbi <= 8'h20;
		14'h1a6f:	ff_dbi <= 8'h20;
		14'h1a70:	ff_dbi <= 8'h20;
		14'h1a71:	ff_dbi <= 8'h20;
		14'h1a72:	ff_dbi <= 8'h20;
		14'h1a73:	ff_dbi <= 8'h20;
		14'h1a74:	ff_dbi <= 8'h20;
		14'h1a75:	ff_dbi <= 8'h20;
		14'h1a76:	ff_dbi <= 8'h20;
		14'h1a77:	ff_dbi <= 8'h20;
		14'h1a78:	ff_dbi <= 8'h20;
		14'h1a79:	ff_dbi <= 8'h20;
		14'h1a7a:	ff_dbi <= 8'h20;
		14'h1a7b:	ff_dbi <= 8'h20;
		14'h1a7c:	ff_dbi <= 8'h20;
		14'h1a7d:	ff_dbi <= 8'h20;
		14'h1a7e:	ff_dbi <= 8'h20;
		14'h1a7f:	ff_dbi <= 8'h20;
		14'h1a80:	ff_dbi <= 8'h20;
		14'h1a81:	ff_dbi <= 8'h20;
		14'h1a82:	ff_dbi <= 8'h20;
		14'h1a83:	ff_dbi <= 8'h20;
		14'h1a84:	ff_dbi <= 8'h20;
		14'h1a85:	ff_dbi <= 8'h20;
		14'h1a86:	ff_dbi <= 8'h20;
		14'h1a87:	ff_dbi <= 8'h20;
		14'h1a88:	ff_dbi <= 8'h20;
		14'h1a89:	ff_dbi <= 8'h20;
		14'h1a8a:	ff_dbi <= 8'h20;
		14'h1a8b:	ff_dbi <= 8'h20;
		14'h1a8c:	ff_dbi <= 8'h20;
		14'h1a8d:	ff_dbi <= 8'h20;
		14'h1a8e:	ff_dbi <= 8'h20;
		14'h1a8f:	ff_dbi <= 8'h20;
		14'h1a90:	ff_dbi <= 8'h20;
		14'h1a91:	ff_dbi <= 8'h20;
		14'h1a92:	ff_dbi <= 8'h20;
		14'h1a93:	ff_dbi <= 8'h20;
		14'h1a94:	ff_dbi <= 8'h20;
		14'h1a95:	ff_dbi <= 8'h20;
		14'h1a96:	ff_dbi <= 8'h20;
		14'h1a97:	ff_dbi <= 8'h20;
		14'h1a98:	ff_dbi <= 8'h20;
		14'h1a99:	ff_dbi <= 8'h20;
		14'h1a9a:	ff_dbi <= 8'h20;
		14'h1a9b:	ff_dbi <= 8'h20;
		14'h1a9c:	ff_dbi <= 8'h20;
		14'h1a9d:	ff_dbi <= 8'h20;
		14'h1a9e:	ff_dbi <= 8'h20;
		14'h1a9f:	ff_dbi <= 8'h20;
		14'h1aa0:	ff_dbi <= 8'h20;
		14'h1aa1:	ff_dbi <= 8'h20;
		14'h1aa2:	ff_dbi <= 8'h20;
		14'h1aa3:	ff_dbi <= 8'h20;
		14'h1aa4:	ff_dbi <= 8'h20;
		14'h1aa5:	ff_dbi <= 8'h20;
		14'h1aa6:	ff_dbi <= 8'h20;
		14'h1aa7:	ff_dbi <= 8'h20;
		14'h1aa8:	ff_dbi <= 8'h20;
		14'h1aa9:	ff_dbi <= 8'h20;
		14'h1aaa:	ff_dbi <= 8'h20;
		14'h1aab:	ff_dbi <= 8'h20;
		14'h1aac:	ff_dbi <= 8'h20;
		14'h1aad:	ff_dbi <= 8'h20;
		14'h1aae:	ff_dbi <= 8'h20;
		14'h1aaf:	ff_dbi <= 8'h20;
		14'h1ab0:	ff_dbi <= 8'h20;
		14'h1ab1:	ff_dbi <= 8'h20;
		14'h1ab2:	ff_dbi <= 8'h20;
		14'h1ab3:	ff_dbi <= 8'h20;
		14'h1ab4:	ff_dbi <= 8'h20;
		14'h1ab5:	ff_dbi <= 8'h20;
		14'h1ab6:	ff_dbi <= 8'h20;
		14'h1ab7:	ff_dbi <= 8'h20;
		14'h1ab8:	ff_dbi <= 8'h20;
		14'h1ab9:	ff_dbi <= 8'h20;
		14'h1aba:	ff_dbi <= 8'h20;
		14'h1abb:	ff_dbi <= 8'h20;
		14'h1abc:	ff_dbi <= 8'h20;
		14'h1abd:	ff_dbi <= 8'h20;
		14'h1abe:	ff_dbi <= 8'h20;
		14'h1abf:	ff_dbi <= 8'h20;
		14'h1ac0:	ff_dbi <= 8'h20;
		14'h1ac1:	ff_dbi <= 8'h20;
		14'h1ac2:	ff_dbi <= 8'h20;
		14'h1ac3:	ff_dbi <= 8'h20;
		14'h1ac4:	ff_dbi <= 8'h20;
		14'h1ac5:	ff_dbi <= 8'h20;
		14'h1ac6:	ff_dbi <= 8'h20;
		14'h1ac7:	ff_dbi <= 8'h20;
		14'h1ac8:	ff_dbi <= 8'h20;
		14'h1ac9:	ff_dbi <= 8'h20;
		14'h1aca:	ff_dbi <= 8'h20;
		14'h1acb:	ff_dbi <= 8'h20;
		14'h1acc:	ff_dbi <= 8'h20;
		14'h1acd:	ff_dbi <= 8'h20;
		14'h1ace:	ff_dbi <= 8'h20;
		14'h1acf:	ff_dbi <= 8'h20;
		14'h1ad0:	ff_dbi <= 8'h20;
		14'h1ad1:	ff_dbi <= 8'h20;
		14'h1ad2:	ff_dbi <= 8'h20;
		14'h1ad3:	ff_dbi <= 8'h20;
		14'h1ad4:	ff_dbi <= 8'h20;
		14'h1ad5:	ff_dbi <= 8'h20;
		14'h1ad6:	ff_dbi <= 8'h20;
		14'h1ad7:	ff_dbi <= 8'h20;
		14'h1ad8:	ff_dbi <= 8'h20;
		14'h1ad9:	ff_dbi <= 8'h20;
		14'h1ada:	ff_dbi <= 8'h20;
		14'h1adb:	ff_dbi <= 8'h20;
		14'h1adc:	ff_dbi <= 8'h20;
		14'h1add:	ff_dbi <= 8'h20;
		14'h1ade:	ff_dbi <= 8'h20;
		14'h1adf:	ff_dbi <= 8'h20;
		14'h1ae0:	ff_dbi <= 8'h20;
		14'h1ae1:	ff_dbi <= 8'h20;
		14'h1ae2:	ff_dbi <= 8'h63;
		14'h1ae3:	ff_dbi <= 8'h6f;
		14'h1ae4:	ff_dbi <= 8'h6c;
		14'h1ae5:	ff_dbi <= 8'h6f;
		14'h1ae6:	ff_dbi <= 8'h72;
		14'h1ae7:	ff_dbi <= 8'h20;
		14'h1ae8:	ff_dbi <= 8'h61;
		14'h1ae9:	ff_dbi <= 8'h75;
		14'h1aea:	ff_dbi <= 8'h74;
		14'h1aeb:	ff_dbi <= 8'h6f;
		14'h1aec:	ff_dbi <= 8'h20;
		14'h1aed:	ff_dbi <= 8'h20;
		14'h1aee:	ff_dbi <= 8'h67;
		14'h1aef:	ff_dbi <= 8'h6f;
		14'h1af0:	ff_dbi <= 8'h74;
		14'h1af1:	ff_dbi <= 8'h6f;
		14'h1af2:	ff_dbi <= 8'h20;
		14'h1af3:	ff_dbi <= 8'h20;
		14'h1af4:	ff_dbi <= 8'h6c;
		14'h1af5:	ff_dbi <= 8'h69;
		14'h1af6:	ff_dbi <= 8'h73;
		14'h1af7:	ff_dbi <= 8'h74;
		14'h1af8:	ff_dbi <= 8'h20;
		14'h1af9:	ff_dbi <= 8'h20;
		14'h1afa:	ff_dbi <= 8'h72;
		14'h1afb:	ff_dbi <= 8'h75;
		14'h1afc:	ff_dbi <= 8'h6e;
		14'h1afd:	ff_dbi <= 8'h20;
		14'h1afe:	ff_dbi <= 8'h20;
		14'h1aff:	ff_dbi <= 8'h20;
		14'h1b00:	ff_dbi <= 8'hd1;
		14'h1b01:	ff_dbi <= 8'h00;
		14'h1b02:	ff_dbi <= 8'h00;
		14'h1b03:	ff_dbi <= 8'h0f;
		14'h1b04:	ff_dbi <= 8'hd1;
		14'h1b05:	ff_dbi <= 8'h00;
		14'h1b06:	ff_dbi <= 8'h01;
		14'h1b07:	ff_dbi <= 8'h0f;
		14'h1b08:	ff_dbi <= 8'hd1;
		14'h1b09:	ff_dbi <= 8'h00;
		14'h1b0a:	ff_dbi <= 8'h02;
		14'h1b0b:	ff_dbi <= 8'h0f;
		14'h1b0c:	ff_dbi <= 8'hd1;
		14'h1b0d:	ff_dbi <= 8'h00;
		14'h1b0e:	ff_dbi <= 8'h03;
		14'h1b0f:	ff_dbi <= 8'h0f;
		14'h1b10:	ff_dbi <= 8'hd1;
		14'h1b11:	ff_dbi <= 8'h00;
		14'h1b12:	ff_dbi <= 8'h04;
		14'h1b13:	ff_dbi <= 8'h0f;
		14'h1b14:	ff_dbi <= 8'hd1;
		14'h1b15:	ff_dbi <= 8'h00;
		14'h1b16:	ff_dbi <= 8'h05;
		14'h1b17:	ff_dbi <= 8'h0f;
		14'h1b18:	ff_dbi <= 8'hd1;
		14'h1b19:	ff_dbi <= 8'h00;
		14'h1b1a:	ff_dbi <= 8'h06;
		14'h1b1b:	ff_dbi <= 8'h0f;
		14'h1b1c:	ff_dbi <= 8'hd1;
		14'h1b1d:	ff_dbi <= 8'h00;
		14'h1b1e:	ff_dbi <= 8'h07;
		14'h1b1f:	ff_dbi <= 8'h0f;
		14'h1b20:	ff_dbi <= 8'hd1;
		14'h1b21:	ff_dbi <= 8'h00;
		14'h1b22:	ff_dbi <= 8'h08;
		14'h1b23:	ff_dbi <= 8'h0f;
		14'h1b24:	ff_dbi <= 8'hd1;
		14'h1b25:	ff_dbi <= 8'h00;
		14'h1b26:	ff_dbi <= 8'h09;
		14'h1b27:	ff_dbi <= 8'h0f;
		14'h1b28:	ff_dbi <= 8'hd1;
		14'h1b29:	ff_dbi <= 8'h00;
		14'h1b2a:	ff_dbi <= 8'h0a;
		14'h1b2b:	ff_dbi <= 8'h0f;
		14'h1b2c:	ff_dbi <= 8'hd1;
		14'h1b2d:	ff_dbi <= 8'h00;
		14'h1b2e:	ff_dbi <= 8'h0b;
		14'h1b2f:	ff_dbi <= 8'h0f;
		14'h1b30:	ff_dbi <= 8'hd1;
		14'h1b31:	ff_dbi <= 8'h00;
		14'h1b32:	ff_dbi <= 8'h0c;
		14'h1b33:	ff_dbi <= 8'h0f;
		14'h1b34:	ff_dbi <= 8'hd1;
		14'h1b35:	ff_dbi <= 8'h00;
		14'h1b36:	ff_dbi <= 8'h0d;
		14'h1b37:	ff_dbi <= 8'h0f;
		14'h1b38:	ff_dbi <= 8'hd1;
		14'h1b39:	ff_dbi <= 8'h00;
		14'h1b3a:	ff_dbi <= 8'h0e;
		14'h1b3b:	ff_dbi <= 8'h0f;
		14'h1b3c:	ff_dbi <= 8'hd1;
		14'h1b3d:	ff_dbi <= 8'h00;
		14'h1b3e:	ff_dbi <= 8'h0f;
		14'h1b3f:	ff_dbi <= 8'h0f;
		14'h1b40:	ff_dbi <= 8'hd1;
		14'h1b41:	ff_dbi <= 8'h00;
		14'h1b42:	ff_dbi <= 8'h10;
		14'h1b43:	ff_dbi <= 8'h0f;
		14'h1b44:	ff_dbi <= 8'hd1;
		14'h1b45:	ff_dbi <= 8'h00;
		14'h1b46:	ff_dbi <= 8'h11;
		14'h1b47:	ff_dbi <= 8'h0f;
		14'h1b48:	ff_dbi <= 8'hd1;
		14'h1b49:	ff_dbi <= 8'h00;
		14'h1b4a:	ff_dbi <= 8'h12;
		14'h1b4b:	ff_dbi <= 8'h0f;
		14'h1b4c:	ff_dbi <= 8'hd1;
		14'h1b4d:	ff_dbi <= 8'h00;
		14'h1b4e:	ff_dbi <= 8'h13;
		14'h1b4f:	ff_dbi <= 8'h0f;
		14'h1b50:	ff_dbi <= 8'hd1;
		14'h1b51:	ff_dbi <= 8'h00;
		14'h1b52:	ff_dbi <= 8'h14;
		14'h1b53:	ff_dbi <= 8'h0f;
		14'h1b54:	ff_dbi <= 8'hd1;
		14'h1b55:	ff_dbi <= 8'h00;
		14'h1b56:	ff_dbi <= 8'h15;
		14'h1b57:	ff_dbi <= 8'h0f;
		14'h1b58:	ff_dbi <= 8'hd1;
		14'h1b59:	ff_dbi <= 8'h00;
		14'h1b5a:	ff_dbi <= 8'h16;
		14'h1b5b:	ff_dbi <= 8'h0f;
		14'h1b5c:	ff_dbi <= 8'hd1;
		14'h1b5d:	ff_dbi <= 8'h00;
		14'h1b5e:	ff_dbi <= 8'h17;
		14'h1b5f:	ff_dbi <= 8'h0f;
		14'h1b60:	ff_dbi <= 8'hd1;
		14'h1b61:	ff_dbi <= 8'h00;
		14'h1b62:	ff_dbi <= 8'h18;
		14'h1b63:	ff_dbi <= 8'h0f;
		14'h1b64:	ff_dbi <= 8'hd1;
		14'h1b65:	ff_dbi <= 8'h00;
		14'h1b66:	ff_dbi <= 8'h19;
		14'h1b67:	ff_dbi <= 8'h0f;
		14'h1b68:	ff_dbi <= 8'hd1;
		14'h1b69:	ff_dbi <= 8'h00;
		14'h1b6a:	ff_dbi <= 8'h1a;
		14'h1b6b:	ff_dbi <= 8'h0f;
		14'h1b6c:	ff_dbi <= 8'hd1;
		14'h1b6d:	ff_dbi <= 8'h00;
		14'h1b6e:	ff_dbi <= 8'h1b;
		14'h1b6f:	ff_dbi <= 8'h0f;
		14'h1b70:	ff_dbi <= 8'hd1;
		14'h1b71:	ff_dbi <= 8'h00;
		14'h1b72:	ff_dbi <= 8'h1c;
		14'h1b73:	ff_dbi <= 8'h0f;
		14'h1b74:	ff_dbi <= 8'hd1;
		14'h1b75:	ff_dbi <= 8'h00;
		14'h1b76:	ff_dbi <= 8'h1d;
		14'h1b77:	ff_dbi <= 8'h0f;
		14'h1b78:	ff_dbi <= 8'hd1;
		14'h1b79:	ff_dbi <= 8'h00;
		14'h1b7a:	ff_dbi <= 8'h1e;
		14'h1b7b:	ff_dbi <= 8'h0f;
		14'h1b7c:	ff_dbi <= 8'hd1;
		14'h1b7d:	ff_dbi <= 8'h00;
		14'h1b7e:	ff_dbi <= 8'h1f;
		14'h1b7f:	ff_dbi <= 8'h0f;
		14'h1b80:	ff_dbi <= 8'h00;
		14'h1b81:	ff_dbi <= 8'h00;
		14'h1b82:	ff_dbi <= 8'h00;
		14'h1b83:	ff_dbi <= 8'h00;
		14'h1b84:	ff_dbi <= 8'h11;
		14'h1b85:	ff_dbi <= 8'h06;
		14'h1b86:	ff_dbi <= 8'h33;
		14'h1b87:	ff_dbi <= 8'h07;
		14'h1b88:	ff_dbi <= 8'h17;
		14'h1b89:	ff_dbi <= 8'h01;
		14'h1b8a:	ff_dbi <= 8'h27;
		14'h1b8b:	ff_dbi <= 8'h03;
		14'h1b8c:	ff_dbi <= 8'h51;
		14'h1b8d:	ff_dbi <= 8'h01;
		14'h1b8e:	ff_dbi <= 8'h27;
		14'h1b8f:	ff_dbi <= 8'h06;
		14'h1b90:	ff_dbi <= 8'h71;
		14'h1b91:	ff_dbi <= 8'h01;
		14'h1b92:	ff_dbi <= 8'h73;
		14'h1b93:	ff_dbi <= 8'h03;
		14'h1b94:	ff_dbi <= 8'h61;
		14'h1b95:	ff_dbi <= 8'h06;
		14'h1b96:	ff_dbi <= 8'h64;
		14'h1b97:	ff_dbi <= 8'h06;
		14'h1b98:	ff_dbi <= 8'h11;
		14'h1b99:	ff_dbi <= 8'h04;
		14'h1b9a:	ff_dbi <= 8'h65;
		14'h1b9b:	ff_dbi <= 8'h02;
		14'h1b9c:	ff_dbi <= 8'h55;
		14'h1b9d:	ff_dbi <= 8'h05;
		14'h1b9e:	ff_dbi <= 8'h77;
		14'h1b9f:	ff_dbi <= 8'h07;
		14'h1ba0:	ff_dbi <= 8'h00;
		14'h1ba1:	ff_dbi <= 8'h00;
		14'h1ba2:	ff_dbi <= 8'h00;
		14'h1ba3:	ff_dbi <= 8'h00;
		14'h1ba4:	ff_dbi <= 8'h00;
		14'h1ba5:	ff_dbi <= 8'h00;
		14'h1ba6:	ff_dbi <= 8'h00;
		14'h1ba7:	ff_dbi <= 8'h00;
		14'h1ba8:	ff_dbi <= 8'h00;
		14'h1ba9:	ff_dbi <= 8'h00;
		14'h1baa:	ff_dbi <= 8'h00;
		14'h1bab:	ff_dbi <= 8'h00;
		14'h1bac:	ff_dbi <= 8'h00;
		14'h1bad:	ff_dbi <= 8'h00;
		14'h1bae:	ff_dbi <= 8'h00;
		14'h1baf:	ff_dbi <= 8'h00;
		14'h1bb0:	ff_dbi <= 8'h00;
		14'h1bb1:	ff_dbi <= 8'h00;
		14'h1bb2:	ff_dbi <= 8'h00;
		14'h1bb3:	ff_dbi <= 8'h00;
		14'h1bb4:	ff_dbi <= 8'h00;
		14'h1bb5:	ff_dbi <= 8'h00;
		14'h1bb6:	ff_dbi <= 8'h00;
		14'h1bb7:	ff_dbi <= 8'h00;
		14'h1bb8:	ff_dbi <= 8'h00;
		14'h1bb9:	ff_dbi <= 8'h00;
		14'h1bba:	ff_dbi <= 8'h00;
		14'h1bbb:	ff_dbi <= 8'h00;
		14'h1bbc:	ff_dbi <= 8'h00;
		14'h1bbd:	ff_dbi <= 8'h00;
		14'h1bbe:	ff_dbi <= 8'h00;
		14'h1bbf:	ff_dbi <= 8'h00;
		14'h1bc0:	ff_dbi <= 8'h00;
		14'h1bc1:	ff_dbi <= 8'h00;
		14'h1bc2:	ff_dbi <= 8'h00;
		14'h1bc3:	ff_dbi <= 8'h00;
		14'h1bc4:	ff_dbi <= 8'h00;
		14'h1bc5:	ff_dbi <= 8'h00;
		14'h1bc6:	ff_dbi <= 8'h00;
		14'h1bc7:	ff_dbi <= 8'h00;
		14'h1bc8:	ff_dbi <= 8'h00;
		14'h1bc9:	ff_dbi <= 8'h00;
		14'h1bca:	ff_dbi <= 8'h00;
		14'h1bcb:	ff_dbi <= 8'h00;
		14'h1bcc:	ff_dbi <= 8'h00;
		14'h1bcd:	ff_dbi <= 8'h00;
		14'h1bce:	ff_dbi <= 8'h00;
		14'h1bcf:	ff_dbi <= 8'h00;
		14'h1bd0:	ff_dbi <= 8'h00;
		14'h1bd1:	ff_dbi <= 8'h00;
		14'h1bd2:	ff_dbi <= 8'h00;
		14'h1bd3:	ff_dbi <= 8'h00;
		14'h1bd4:	ff_dbi <= 8'h00;
		14'h1bd5:	ff_dbi <= 8'h00;
		14'h1bd6:	ff_dbi <= 8'h00;
		14'h1bd7:	ff_dbi <= 8'h00;
		14'h1bd8:	ff_dbi <= 8'h00;
		14'h1bd9:	ff_dbi <= 8'h00;
		14'h1bda:	ff_dbi <= 8'h00;
		14'h1bdb:	ff_dbi <= 8'h00;
		14'h1bdc:	ff_dbi <= 8'h00;
		14'h1bdd:	ff_dbi <= 8'h00;
		14'h1bde:	ff_dbi <= 8'h00;
		14'h1bdf:	ff_dbi <= 8'h00;
		14'h1be0:	ff_dbi <= 8'h00;
		14'h1be1:	ff_dbi <= 8'h00;
		14'h1be2:	ff_dbi <= 8'h00;
		14'h1be3:	ff_dbi <= 8'h00;
		14'h1be4:	ff_dbi <= 8'h00;
		14'h1be5:	ff_dbi <= 8'h00;
		14'h1be6:	ff_dbi <= 8'h00;
		14'h1be7:	ff_dbi <= 8'h00;
		14'h1be8:	ff_dbi <= 8'h00;
		14'h1be9:	ff_dbi <= 8'h00;
		14'h1bea:	ff_dbi <= 8'h00;
		14'h1beb:	ff_dbi <= 8'h00;
		14'h1bec:	ff_dbi <= 8'h00;
		14'h1bed:	ff_dbi <= 8'h00;
		14'h1bee:	ff_dbi <= 8'h00;
		14'h1bef:	ff_dbi <= 8'h00;
		14'h1bf0:	ff_dbi <= 8'h00;
		14'h1bf1:	ff_dbi <= 8'h00;
		14'h1bf2:	ff_dbi <= 8'h00;
		14'h1bf3:	ff_dbi <= 8'h00;
		14'h1bf4:	ff_dbi <= 8'h00;
		14'h1bf5:	ff_dbi <= 8'h00;
		14'h1bf6:	ff_dbi <= 8'h00;
		14'h1bf7:	ff_dbi <= 8'h00;
		14'h1bf8:	ff_dbi <= 8'h00;
		14'h1bf9:	ff_dbi <= 8'h00;
		14'h1bfa:	ff_dbi <= 8'h00;
		14'h1bfb:	ff_dbi <= 8'h00;
		14'h1bfc:	ff_dbi <= 8'h00;
		14'h1bfd:	ff_dbi <= 8'h00;
		14'h1bfe:	ff_dbi <= 8'h00;
		14'h1bff:	ff_dbi <= 8'h00;
		14'h1c00:	ff_dbi <= 8'h00;
		14'h1c01:	ff_dbi <= 8'h00;
		14'h1c02:	ff_dbi <= 8'h00;
		14'h1c03:	ff_dbi <= 8'h00;
		14'h1c04:	ff_dbi <= 8'h00;
		14'h1c05:	ff_dbi <= 8'h00;
		14'h1c06:	ff_dbi <= 8'h00;
		14'h1c07:	ff_dbi <= 8'h00;
		14'h1c08:	ff_dbi <= 8'h00;
		14'h1c09:	ff_dbi <= 8'h00;
		14'h1c0a:	ff_dbi <= 8'h00;
		14'h1c0b:	ff_dbi <= 8'h00;
		14'h1c0c:	ff_dbi <= 8'h00;
		14'h1c0d:	ff_dbi <= 8'h00;
		14'h1c0e:	ff_dbi <= 8'h00;
		14'h1c0f:	ff_dbi <= 8'h00;
		14'h1c10:	ff_dbi <= 8'h00;
		14'h1c11:	ff_dbi <= 8'h00;
		14'h1c12:	ff_dbi <= 8'h00;
		14'h1c13:	ff_dbi <= 8'h00;
		14'h1c14:	ff_dbi <= 8'h00;
		14'h1c15:	ff_dbi <= 8'h00;
		14'h1c16:	ff_dbi <= 8'h00;
		14'h1c17:	ff_dbi <= 8'h00;
		14'h1c18:	ff_dbi <= 8'h00;
		14'h1c19:	ff_dbi <= 8'h00;
		14'h1c1a:	ff_dbi <= 8'h00;
		14'h1c1b:	ff_dbi <= 8'h00;
		14'h1c1c:	ff_dbi <= 8'h00;
		14'h1c1d:	ff_dbi <= 8'h00;
		14'h1c1e:	ff_dbi <= 8'h00;
		14'h1c1f:	ff_dbi <= 8'h00;
		14'h1c20:	ff_dbi <= 8'h00;
		14'h1c21:	ff_dbi <= 8'h00;
		14'h1c22:	ff_dbi <= 8'h00;
		14'h1c23:	ff_dbi <= 8'h00;
		14'h1c24:	ff_dbi <= 8'h00;
		14'h1c25:	ff_dbi <= 8'h00;
		14'h1c26:	ff_dbi <= 8'h00;
		14'h1c27:	ff_dbi <= 8'h00;
		14'h1c28:	ff_dbi <= 8'h00;
		14'h1c29:	ff_dbi <= 8'h00;
		14'h1c2a:	ff_dbi <= 8'h00;
		14'h1c2b:	ff_dbi <= 8'h00;
		14'h1c2c:	ff_dbi <= 8'h00;
		14'h1c2d:	ff_dbi <= 8'h00;
		14'h1c2e:	ff_dbi <= 8'h00;
		14'h1c2f:	ff_dbi <= 8'h00;
		14'h1c30:	ff_dbi <= 8'h00;
		14'h1c31:	ff_dbi <= 8'h00;
		14'h1c32:	ff_dbi <= 8'h00;
		14'h1c33:	ff_dbi <= 8'h00;
		14'h1c34:	ff_dbi <= 8'h00;
		14'h1c35:	ff_dbi <= 8'h00;
		14'h1c36:	ff_dbi <= 8'h00;
		14'h1c37:	ff_dbi <= 8'h00;
		14'h1c38:	ff_dbi <= 8'h00;
		14'h1c39:	ff_dbi <= 8'h00;
		14'h1c3a:	ff_dbi <= 8'h00;
		14'h1c3b:	ff_dbi <= 8'h00;
		14'h1c3c:	ff_dbi <= 8'h00;
		14'h1c3d:	ff_dbi <= 8'h00;
		14'h1c3e:	ff_dbi <= 8'h00;
		14'h1c3f:	ff_dbi <= 8'h00;
		14'h1c40:	ff_dbi <= 8'h00;
		14'h1c41:	ff_dbi <= 8'h00;
		14'h1c42:	ff_dbi <= 8'h00;
		14'h1c43:	ff_dbi <= 8'h00;
		14'h1c44:	ff_dbi <= 8'h00;
		14'h1c45:	ff_dbi <= 8'h00;
		14'h1c46:	ff_dbi <= 8'h00;
		14'h1c47:	ff_dbi <= 8'h00;
		14'h1c48:	ff_dbi <= 8'h00;
		14'h1c49:	ff_dbi <= 8'h00;
		14'h1c4a:	ff_dbi <= 8'h00;
		14'h1c4b:	ff_dbi <= 8'h00;
		14'h1c4c:	ff_dbi <= 8'h00;
		14'h1c4d:	ff_dbi <= 8'h00;
		14'h1c4e:	ff_dbi <= 8'h00;
		14'h1c4f:	ff_dbi <= 8'h00;
		14'h1c50:	ff_dbi <= 8'h00;
		14'h1c51:	ff_dbi <= 8'h00;
		14'h1c52:	ff_dbi <= 8'h00;
		14'h1c53:	ff_dbi <= 8'h00;
		14'h1c54:	ff_dbi <= 8'h00;
		14'h1c55:	ff_dbi <= 8'h00;
		14'h1c56:	ff_dbi <= 8'h00;
		14'h1c57:	ff_dbi <= 8'h00;
		14'h1c58:	ff_dbi <= 8'h00;
		14'h1c59:	ff_dbi <= 8'h00;
		14'h1c5a:	ff_dbi <= 8'h00;
		14'h1c5b:	ff_dbi <= 8'h00;
		14'h1c5c:	ff_dbi <= 8'h00;
		14'h1c5d:	ff_dbi <= 8'h00;
		14'h1c5e:	ff_dbi <= 8'h00;
		14'h1c5f:	ff_dbi <= 8'h00;
		14'h1c60:	ff_dbi <= 8'h00;
		14'h1c61:	ff_dbi <= 8'h00;
		14'h1c62:	ff_dbi <= 8'h00;
		14'h1c63:	ff_dbi <= 8'h00;
		14'h1c64:	ff_dbi <= 8'h00;
		14'h1c65:	ff_dbi <= 8'h00;
		14'h1c66:	ff_dbi <= 8'h00;
		14'h1c67:	ff_dbi <= 8'h00;
		14'h1c68:	ff_dbi <= 8'h00;
		14'h1c69:	ff_dbi <= 8'h00;
		14'h1c6a:	ff_dbi <= 8'h00;
		14'h1c6b:	ff_dbi <= 8'h00;
		14'h1c6c:	ff_dbi <= 8'h00;
		14'h1c6d:	ff_dbi <= 8'h00;
		14'h1c6e:	ff_dbi <= 8'h00;
		14'h1c6f:	ff_dbi <= 8'h00;
		14'h1c70:	ff_dbi <= 8'h00;
		14'h1c71:	ff_dbi <= 8'h00;
		14'h1c72:	ff_dbi <= 8'h00;
		14'h1c73:	ff_dbi <= 8'h00;
		14'h1c74:	ff_dbi <= 8'h00;
		14'h1c75:	ff_dbi <= 8'h00;
		14'h1c76:	ff_dbi <= 8'h00;
		14'h1c77:	ff_dbi <= 8'h00;
		14'h1c78:	ff_dbi <= 8'h00;
		14'h1c79:	ff_dbi <= 8'h00;
		14'h1c7a:	ff_dbi <= 8'h00;
		14'h1c7b:	ff_dbi <= 8'h00;
		14'h1c7c:	ff_dbi <= 8'h00;
		14'h1c7d:	ff_dbi <= 8'h00;
		14'h1c7e:	ff_dbi <= 8'h00;
		14'h1c7f:	ff_dbi <= 8'h00;
		14'h1c80:	ff_dbi <= 8'h00;
		14'h1c81:	ff_dbi <= 8'h00;
		14'h1c82:	ff_dbi <= 8'h00;
		14'h1c83:	ff_dbi <= 8'h00;
		14'h1c84:	ff_dbi <= 8'h00;
		14'h1c85:	ff_dbi <= 8'h00;
		14'h1c86:	ff_dbi <= 8'h00;
		14'h1c87:	ff_dbi <= 8'h00;
		14'h1c88:	ff_dbi <= 8'h00;
		14'h1c89:	ff_dbi <= 8'h00;
		14'h1c8a:	ff_dbi <= 8'h00;
		14'h1c8b:	ff_dbi <= 8'h00;
		14'h1c8c:	ff_dbi <= 8'h00;
		14'h1c8d:	ff_dbi <= 8'h00;
		14'h1c8e:	ff_dbi <= 8'h00;
		14'h1c8f:	ff_dbi <= 8'h00;
		14'h1c90:	ff_dbi <= 8'h00;
		14'h1c91:	ff_dbi <= 8'h00;
		14'h1c92:	ff_dbi <= 8'h00;
		14'h1c93:	ff_dbi <= 8'h00;
		14'h1c94:	ff_dbi <= 8'h00;
		14'h1c95:	ff_dbi <= 8'h00;
		14'h1c96:	ff_dbi <= 8'h00;
		14'h1c97:	ff_dbi <= 8'h00;
		14'h1c98:	ff_dbi <= 8'h00;
		14'h1c99:	ff_dbi <= 8'h00;
		14'h1c9a:	ff_dbi <= 8'h00;
		14'h1c9b:	ff_dbi <= 8'h00;
		14'h1c9c:	ff_dbi <= 8'h00;
		14'h1c9d:	ff_dbi <= 8'h00;
		14'h1c9e:	ff_dbi <= 8'h00;
		14'h1c9f:	ff_dbi <= 8'h00;
		14'h1ca0:	ff_dbi <= 8'h00;
		14'h1ca1:	ff_dbi <= 8'h00;
		14'h1ca2:	ff_dbi <= 8'h00;
		14'h1ca3:	ff_dbi <= 8'h00;
		14'h1ca4:	ff_dbi <= 8'h00;
		14'h1ca5:	ff_dbi <= 8'h00;
		14'h1ca6:	ff_dbi <= 8'h00;
		14'h1ca7:	ff_dbi <= 8'h00;
		14'h1ca8:	ff_dbi <= 8'h00;
		14'h1ca9:	ff_dbi <= 8'h00;
		14'h1caa:	ff_dbi <= 8'h00;
		14'h1cab:	ff_dbi <= 8'h00;
		14'h1cac:	ff_dbi <= 8'h00;
		14'h1cad:	ff_dbi <= 8'h00;
		14'h1cae:	ff_dbi <= 8'h00;
		14'h1caf:	ff_dbi <= 8'h00;
		14'h1cb0:	ff_dbi <= 8'h00;
		14'h1cb1:	ff_dbi <= 8'h00;
		14'h1cb2:	ff_dbi <= 8'h00;
		14'h1cb3:	ff_dbi <= 8'h00;
		14'h1cb4:	ff_dbi <= 8'h00;
		14'h1cb5:	ff_dbi <= 8'h00;
		14'h1cb6:	ff_dbi <= 8'h00;
		14'h1cb7:	ff_dbi <= 8'h00;
		14'h1cb8:	ff_dbi <= 8'h00;
		14'h1cb9:	ff_dbi <= 8'h00;
		14'h1cba:	ff_dbi <= 8'h00;
		14'h1cbb:	ff_dbi <= 8'h00;
		14'h1cbc:	ff_dbi <= 8'h00;
		14'h1cbd:	ff_dbi <= 8'h00;
		14'h1cbe:	ff_dbi <= 8'h00;
		14'h1cbf:	ff_dbi <= 8'h00;
		14'h1cc0:	ff_dbi <= 8'h00;
		14'h1cc1:	ff_dbi <= 8'h00;
		14'h1cc2:	ff_dbi <= 8'h00;
		14'h1cc3:	ff_dbi <= 8'h00;
		14'h1cc4:	ff_dbi <= 8'h00;
		14'h1cc5:	ff_dbi <= 8'h00;
		14'h1cc6:	ff_dbi <= 8'h00;
		14'h1cc7:	ff_dbi <= 8'h00;
		14'h1cc8:	ff_dbi <= 8'h00;
		14'h1cc9:	ff_dbi <= 8'h00;
		14'h1cca:	ff_dbi <= 8'h00;
		14'h1ccb:	ff_dbi <= 8'h00;
		14'h1ccc:	ff_dbi <= 8'h00;
		14'h1ccd:	ff_dbi <= 8'h00;
		14'h1cce:	ff_dbi <= 8'h00;
		14'h1ccf:	ff_dbi <= 8'h00;
		14'h1cd0:	ff_dbi <= 8'h00;
		14'h1cd1:	ff_dbi <= 8'h00;
		14'h1cd2:	ff_dbi <= 8'h00;
		14'h1cd3:	ff_dbi <= 8'h00;
		14'h1cd4:	ff_dbi <= 8'h00;
		14'h1cd5:	ff_dbi <= 8'h00;
		14'h1cd6:	ff_dbi <= 8'h00;
		14'h1cd7:	ff_dbi <= 8'h00;
		14'h1cd8:	ff_dbi <= 8'h00;
		14'h1cd9:	ff_dbi <= 8'h00;
		14'h1cda:	ff_dbi <= 8'h00;
		14'h1cdb:	ff_dbi <= 8'h00;
		14'h1cdc:	ff_dbi <= 8'h00;
		14'h1cdd:	ff_dbi <= 8'h00;
		14'h1cde:	ff_dbi <= 8'h00;
		14'h1cdf:	ff_dbi <= 8'h00;
		14'h1ce0:	ff_dbi <= 8'h00;
		14'h1ce1:	ff_dbi <= 8'h00;
		14'h1ce2:	ff_dbi <= 8'h00;
		14'h1ce3:	ff_dbi <= 8'h00;
		14'h1ce4:	ff_dbi <= 8'h00;
		14'h1ce5:	ff_dbi <= 8'h00;
		14'h1ce6:	ff_dbi <= 8'h00;
		14'h1ce7:	ff_dbi <= 8'h00;
		14'h1ce8:	ff_dbi <= 8'h00;
		14'h1ce9:	ff_dbi <= 8'h00;
		14'h1cea:	ff_dbi <= 8'h00;
		14'h1ceb:	ff_dbi <= 8'h00;
		14'h1cec:	ff_dbi <= 8'h00;
		14'h1ced:	ff_dbi <= 8'h00;
		14'h1cee:	ff_dbi <= 8'h00;
		14'h1cef:	ff_dbi <= 8'h00;
		14'h1cf0:	ff_dbi <= 8'h00;
		14'h1cf1:	ff_dbi <= 8'h00;
		14'h1cf2:	ff_dbi <= 8'h00;
		14'h1cf3:	ff_dbi <= 8'h00;
		14'h1cf4:	ff_dbi <= 8'h00;
		14'h1cf5:	ff_dbi <= 8'h00;
		14'h1cf6:	ff_dbi <= 8'h00;
		14'h1cf7:	ff_dbi <= 8'h00;
		14'h1cf8:	ff_dbi <= 8'h00;
		14'h1cf9:	ff_dbi <= 8'h00;
		14'h1cfa:	ff_dbi <= 8'h00;
		14'h1cfb:	ff_dbi <= 8'h00;
		14'h1cfc:	ff_dbi <= 8'h00;
		14'h1cfd:	ff_dbi <= 8'h00;
		14'h1cfe:	ff_dbi <= 8'h00;
		14'h1cff:	ff_dbi <= 8'h00;
		14'h1d00:	ff_dbi <= 8'h00;
		14'h1d01:	ff_dbi <= 8'h00;
		14'h1d02:	ff_dbi <= 8'h00;
		14'h1d03:	ff_dbi <= 8'h00;
		14'h1d04:	ff_dbi <= 8'h00;
		14'h1d05:	ff_dbi <= 8'h00;
		14'h1d06:	ff_dbi <= 8'h00;
		14'h1d07:	ff_dbi <= 8'h00;
		14'h1d08:	ff_dbi <= 8'h00;
		14'h1d09:	ff_dbi <= 8'h00;
		14'h1d0a:	ff_dbi <= 8'h00;
		14'h1d0b:	ff_dbi <= 8'h00;
		14'h1d0c:	ff_dbi <= 8'h00;
		14'h1d0d:	ff_dbi <= 8'h00;
		14'h1d0e:	ff_dbi <= 8'h00;
		14'h1d0f:	ff_dbi <= 8'h00;
		14'h1d10:	ff_dbi <= 8'h00;
		14'h1d11:	ff_dbi <= 8'h00;
		14'h1d12:	ff_dbi <= 8'h00;
		14'h1d13:	ff_dbi <= 8'h00;
		14'h1d14:	ff_dbi <= 8'h00;
		14'h1d15:	ff_dbi <= 8'h00;
		14'h1d16:	ff_dbi <= 8'h00;
		14'h1d17:	ff_dbi <= 8'h00;
		14'h1d18:	ff_dbi <= 8'h00;
		14'h1d19:	ff_dbi <= 8'h00;
		14'h1d1a:	ff_dbi <= 8'h00;
		14'h1d1b:	ff_dbi <= 8'h00;
		14'h1d1c:	ff_dbi <= 8'h00;
		14'h1d1d:	ff_dbi <= 8'h00;
		14'h1d1e:	ff_dbi <= 8'h00;
		14'h1d1f:	ff_dbi <= 8'h00;
		14'h1d20:	ff_dbi <= 8'h00;
		14'h1d21:	ff_dbi <= 8'h00;
		14'h1d22:	ff_dbi <= 8'h00;
		14'h1d23:	ff_dbi <= 8'h00;
		14'h1d24:	ff_dbi <= 8'h00;
		14'h1d25:	ff_dbi <= 8'h00;
		14'h1d26:	ff_dbi <= 8'h00;
		14'h1d27:	ff_dbi <= 8'h00;
		14'h1d28:	ff_dbi <= 8'h00;
		14'h1d29:	ff_dbi <= 8'h00;
		14'h1d2a:	ff_dbi <= 8'h00;
		14'h1d2b:	ff_dbi <= 8'h00;
		14'h1d2c:	ff_dbi <= 8'h00;
		14'h1d2d:	ff_dbi <= 8'h00;
		14'h1d2e:	ff_dbi <= 8'h00;
		14'h1d2f:	ff_dbi <= 8'h00;
		14'h1d30:	ff_dbi <= 8'h00;
		14'h1d31:	ff_dbi <= 8'h00;
		14'h1d32:	ff_dbi <= 8'h00;
		14'h1d33:	ff_dbi <= 8'h00;
		14'h1d34:	ff_dbi <= 8'h00;
		14'h1d35:	ff_dbi <= 8'h00;
		14'h1d36:	ff_dbi <= 8'h00;
		14'h1d37:	ff_dbi <= 8'h00;
		14'h1d38:	ff_dbi <= 8'h00;
		14'h1d39:	ff_dbi <= 8'h00;
		14'h1d3a:	ff_dbi <= 8'h00;
		14'h1d3b:	ff_dbi <= 8'h00;
		14'h1d3c:	ff_dbi <= 8'h00;
		14'h1d3d:	ff_dbi <= 8'h00;
		14'h1d3e:	ff_dbi <= 8'h00;
		14'h1d3f:	ff_dbi <= 8'h00;
		14'h1d40:	ff_dbi <= 8'h00;
		14'h1d41:	ff_dbi <= 8'h00;
		14'h1d42:	ff_dbi <= 8'h00;
		14'h1d43:	ff_dbi <= 8'h00;
		14'h1d44:	ff_dbi <= 8'h00;
		14'h1d45:	ff_dbi <= 8'h00;
		14'h1d46:	ff_dbi <= 8'h00;
		14'h1d47:	ff_dbi <= 8'h00;
		14'h1d48:	ff_dbi <= 8'h00;
		14'h1d49:	ff_dbi <= 8'h00;
		14'h1d4a:	ff_dbi <= 8'h00;
		14'h1d4b:	ff_dbi <= 8'h00;
		14'h1d4c:	ff_dbi <= 8'h00;
		14'h1d4d:	ff_dbi <= 8'h00;
		14'h1d4e:	ff_dbi <= 8'h00;
		14'h1d4f:	ff_dbi <= 8'h00;
		14'h1d50:	ff_dbi <= 8'h00;
		14'h1d51:	ff_dbi <= 8'h00;
		14'h1d52:	ff_dbi <= 8'h00;
		14'h1d53:	ff_dbi <= 8'h00;
		14'h1d54:	ff_dbi <= 8'h00;
		14'h1d55:	ff_dbi <= 8'h00;
		14'h1d56:	ff_dbi <= 8'h00;
		14'h1d57:	ff_dbi <= 8'h00;
		14'h1d58:	ff_dbi <= 8'h00;
		14'h1d59:	ff_dbi <= 8'h00;
		14'h1d5a:	ff_dbi <= 8'h00;
		14'h1d5b:	ff_dbi <= 8'h00;
		14'h1d5c:	ff_dbi <= 8'h00;
		14'h1d5d:	ff_dbi <= 8'h00;
		14'h1d5e:	ff_dbi <= 8'h00;
		14'h1d5f:	ff_dbi <= 8'h00;
		14'h1d60:	ff_dbi <= 8'h00;
		14'h1d61:	ff_dbi <= 8'h00;
		14'h1d62:	ff_dbi <= 8'h00;
		14'h1d63:	ff_dbi <= 8'h00;
		14'h1d64:	ff_dbi <= 8'h00;
		14'h1d65:	ff_dbi <= 8'h00;
		14'h1d66:	ff_dbi <= 8'h00;
		14'h1d67:	ff_dbi <= 8'h00;
		14'h1d68:	ff_dbi <= 8'h00;
		14'h1d69:	ff_dbi <= 8'h00;
		14'h1d6a:	ff_dbi <= 8'h00;
		14'h1d6b:	ff_dbi <= 8'h00;
		14'h1d6c:	ff_dbi <= 8'h00;
		14'h1d6d:	ff_dbi <= 8'h00;
		14'h1d6e:	ff_dbi <= 8'h00;
		14'h1d6f:	ff_dbi <= 8'h00;
		14'h1d70:	ff_dbi <= 8'h00;
		14'h1d71:	ff_dbi <= 8'h00;
		14'h1d72:	ff_dbi <= 8'h00;
		14'h1d73:	ff_dbi <= 8'h00;
		14'h1d74:	ff_dbi <= 8'h00;
		14'h1d75:	ff_dbi <= 8'h00;
		14'h1d76:	ff_dbi <= 8'h00;
		14'h1d77:	ff_dbi <= 8'h00;
		14'h1d78:	ff_dbi <= 8'h00;
		14'h1d79:	ff_dbi <= 8'h00;
		14'h1d7a:	ff_dbi <= 8'h00;
		14'h1d7b:	ff_dbi <= 8'h00;
		14'h1d7c:	ff_dbi <= 8'h00;
		14'h1d7d:	ff_dbi <= 8'h00;
		14'h1d7e:	ff_dbi <= 8'h00;
		14'h1d7f:	ff_dbi <= 8'h00;
		14'h1d80:	ff_dbi <= 8'h00;
		14'h1d81:	ff_dbi <= 8'h00;
		14'h1d82:	ff_dbi <= 8'h00;
		14'h1d83:	ff_dbi <= 8'h00;
		14'h1d84:	ff_dbi <= 8'h00;
		14'h1d85:	ff_dbi <= 8'h00;
		14'h1d86:	ff_dbi <= 8'h00;
		14'h1d87:	ff_dbi <= 8'h00;
		14'h1d88:	ff_dbi <= 8'h00;
		14'h1d89:	ff_dbi <= 8'h00;
		14'h1d8a:	ff_dbi <= 8'h00;
		14'h1d8b:	ff_dbi <= 8'h00;
		14'h1d8c:	ff_dbi <= 8'h00;
		14'h1d8d:	ff_dbi <= 8'h00;
		14'h1d8e:	ff_dbi <= 8'h00;
		14'h1d8f:	ff_dbi <= 8'h00;
		14'h1d90:	ff_dbi <= 8'h00;
		14'h1d91:	ff_dbi <= 8'h00;
		14'h1d92:	ff_dbi <= 8'h00;
		14'h1d93:	ff_dbi <= 8'h00;
		14'h1d94:	ff_dbi <= 8'h00;
		14'h1d95:	ff_dbi <= 8'h00;
		14'h1d96:	ff_dbi <= 8'h00;
		14'h1d97:	ff_dbi <= 8'h00;
		14'h1d98:	ff_dbi <= 8'h00;
		14'h1d99:	ff_dbi <= 8'h00;
		14'h1d9a:	ff_dbi <= 8'h00;
		14'h1d9b:	ff_dbi <= 8'h00;
		14'h1d9c:	ff_dbi <= 8'h00;
		14'h1d9d:	ff_dbi <= 8'h00;
		14'h1d9e:	ff_dbi <= 8'h00;
		14'h1d9f:	ff_dbi <= 8'h00;
		14'h1da0:	ff_dbi <= 8'h00;
		14'h1da1:	ff_dbi <= 8'h00;
		14'h1da2:	ff_dbi <= 8'h00;
		14'h1da3:	ff_dbi <= 8'h00;
		14'h1da4:	ff_dbi <= 8'h00;
		14'h1da5:	ff_dbi <= 8'h00;
		14'h1da6:	ff_dbi <= 8'h00;
		14'h1da7:	ff_dbi <= 8'h00;
		14'h1da8:	ff_dbi <= 8'h00;
		14'h1da9:	ff_dbi <= 8'h00;
		14'h1daa:	ff_dbi <= 8'h00;
		14'h1dab:	ff_dbi <= 8'h00;
		14'h1dac:	ff_dbi <= 8'h00;
		14'h1dad:	ff_dbi <= 8'h00;
		14'h1dae:	ff_dbi <= 8'h00;
		14'h1daf:	ff_dbi <= 8'h00;
		14'h1db0:	ff_dbi <= 8'h00;
		14'h1db1:	ff_dbi <= 8'h00;
		14'h1db2:	ff_dbi <= 8'h00;
		14'h1db3:	ff_dbi <= 8'h00;
		14'h1db4:	ff_dbi <= 8'h00;
		14'h1db5:	ff_dbi <= 8'h00;
		14'h1db6:	ff_dbi <= 8'h00;
		14'h1db7:	ff_dbi <= 8'h00;
		14'h1db8:	ff_dbi <= 8'h00;
		14'h1db9:	ff_dbi <= 8'h00;
		14'h1dba:	ff_dbi <= 8'h00;
		14'h1dbb:	ff_dbi <= 8'h00;
		14'h1dbc:	ff_dbi <= 8'h00;
		14'h1dbd:	ff_dbi <= 8'h00;
		14'h1dbe:	ff_dbi <= 8'h00;
		14'h1dbf:	ff_dbi <= 8'h00;
		14'h1dc0:	ff_dbi <= 8'h00;
		14'h1dc1:	ff_dbi <= 8'h00;
		14'h1dc2:	ff_dbi <= 8'h00;
		14'h1dc3:	ff_dbi <= 8'h00;
		14'h1dc4:	ff_dbi <= 8'h00;
		14'h1dc5:	ff_dbi <= 8'h00;
		14'h1dc6:	ff_dbi <= 8'h00;
		14'h1dc7:	ff_dbi <= 8'h00;
		14'h1dc8:	ff_dbi <= 8'h00;
		14'h1dc9:	ff_dbi <= 8'h00;
		14'h1dca:	ff_dbi <= 8'h00;
		14'h1dcb:	ff_dbi <= 8'h00;
		14'h1dcc:	ff_dbi <= 8'h00;
		14'h1dcd:	ff_dbi <= 8'h00;
		14'h1dce:	ff_dbi <= 8'h00;
		14'h1dcf:	ff_dbi <= 8'h00;
		14'h1dd0:	ff_dbi <= 8'h00;
		14'h1dd1:	ff_dbi <= 8'h00;
		14'h1dd2:	ff_dbi <= 8'h00;
		14'h1dd3:	ff_dbi <= 8'h00;
		14'h1dd4:	ff_dbi <= 8'h00;
		14'h1dd5:	ff_dbi <= 8'h00;
		14'h1dd6:	ff_dbi <= 8'h00;
		14'h1dd7:	ff_dbi <= 8'h00;
		14'h1dd8:	ff_dbi <= 8'h00;
		14'h1dd9:	ff_dbi <= 8'h00;
		14'h1dda:	ff_dbi <= 8'h00;
		14'h1ddb:	ff_dbi <= 8'h00;
		14'h1ddc:	ff_dbi <= 8'h00;
		14'h1ddd:	ff_dbi <= 8'h00;
		14'h1dde:	ff_dbi <= 8'h00;
		14'h1ddf:	ff_dbi <= 8'h00;
		14'h1de0:	ff_dbi <= 8'h00;
		14'h1de1:	ff_dbi <= 8'h00;
		14'h1de2:	ff_dbi <= 8'h00;
		14'h1de3:	ff_dbi <= 8'h00;
		14'h1de4:	ff_dbi <= 8'h00;
		14'h1de5:	ff_dbi <= 8'h00;
		14'h1de6:	ff_dbi <= 8'h00;
		14'h1de7:	ff_dbi <= 8'h00;
		14'h1de8:	ff_dbi <= 8'h00;
		14'h1de9:	ff_dbi <= 8'h00;
		14'h1dea:	ff_dbi <= 8'h00;
		14'h1deb:	ff_dbi <= 8'h00;
		14'h1dec:	ff_dbi <= 8'h00;
		14'h1ded:	ff_dbi <= 8'h00;
		14'h1dee:	ff_dbi <= 8'h00;
		14'h1def:	ff_dbi <= 8'h00;
		14'h1df0:	ff_dbi <= 8'h00;
		14'h1df1:	ff_dbi <= 8'h00;
		14'h1df2:	ff_dbi <= 8'h00;
		14'h1df3:	ff_dbi <= 8'h00;
		14'h1df4:	ff_dbi <= 8'h00;
		14'h1df5:	ff_dbi <= 8'h00;
		14'h1df6:	ff_dbi <= 8'h00;
		14'h1df7:	ff_dbi <= 8'h00;
		14'h1df8:	ff_dbi <= 8'h00;
		14'h1df9:	ff_dbi <= 8'h00;
		14'h1dfa:	ff_dbi <= 8'h00;
		14'h1dfb:	ff_dbi <= 8'h00;
		14'h1dfc:	ff_dbi <= 8'h00;
		14'h1dfd:	ff_dbi <= 8'h00;
		14'h1dfe:	ff_dbi <= 8'h00;
		14'h1dff:	ff_dbi <= 8'h00;
		14'h1e00:	ff_dbi <= 8'h00;
		14'h1e01:	ff_dbi <= 8'h00;
		14'h1e02:	ff_dbi <= 8'h00;
		14'h1e03:	ff_dbi <= 8'h00;
		14'h1e04:	ff_dbi <= 8'h00;
		14'h1e05:	ff_dbi <= 8'h00;
		14'h1e06:	ff_dbi <= 8'h00;
		14'h1e07:	ff_dbi <= 8'h00;
		14'h1e08:	ff_dbi <= 8'h00;
		14'h1e09:	ff_dbi <= 8'h00;
		14'h1e0a:	ff_dbi <= 8'h00;
		14'h1e0b:	ff_dbi <= 8'h00;
		14'h1e0c:	ff_dbi <= 8'h00;
		14'h1e0d:	ff_dbi <= 8'h00;
		14'h1e0e:	ff_dbi <= 8'h00;
		14'h1e0f:	ff_dbi <= 8'h00;
		14'h1e10:	ff_dbi <= 8'h00;
		14'h1e11:	ff_dbi <= 8'h00;
		14'h1e12:	ff_dbi <= 8'h00;
		14'h1e13:	ff_dbi <= 8'h00;
		14'h1e14:	ff_dbi <= 8'h00;
		14'h1e15:	ff_dbi <= 8'h00;
		14'h1e16:	ff_dbi <= 8'h00;
		14'h1e17:	ff_dbi <= 8'h00;
		14'h1e18:	ff_dbi <= 8'h00;
		14'h1e19:	ff_dbi <= 8'h00;
		14'h1e1a:	ff_dbi <= 8'h00;
		14'h1e1b:	ff_dbi <= 8'h00;
		14'h1e1c:	ff_dbi <= 8'h00;
		14'h1e1d:	ff_dbi <= 8'h00;
		14'h1e1e:	ff_dbi <= 8'h00;
		14'h1e1f:	ff_dbi <= 8'h00;
		14'h1e20:	ff_dbi <= 8'h00;
		14'h1e21:	ff_dbi <= 8'h00;
		14'h1e22:	ff_dbi <= 8'h00;
		14'h1e23:	ff_dbi <= 8'h00;
		14'h1e24:	ff_dbi <= 8'h00;
		14'h1e25:	ff_dbi <= 8'h00;
		14'h1e26:	ff_dbi <= 8'h00;
		14'h1e27:	ff_dbi <= 8'h00;
		14'h1e28:	ff_dbi <= 8'h00;
		14'h1e29:	ff_dbi <= 8'h00;
		14'h1e2a:	ff_dbi <= 8'h00;
		14'h1e2b:	ff_dbi <= 8'h00;
		14'h1e2c:	ff_dbi <= 8'h00;
		14'h1e2d:	ff_dbi <= 8'h00;
		14'h1e2e:	ff_dbi <= 8'h00;
		14'h1e2f:	ff_dbi <= 8'h00;
		14'h1e30:	ff_dbi <= 8'h00;
		14'h1e31:	ff_dbi <= 8'h00;
		14'h1e32:	ff_dbi <= 8'h00;
		14'h1e33:	ff_dbi <= 8'h00;
		14'h1e34:	ff_dbi <= 8'h00;
		14'h1e35:	ff_dbi <= 8'h00;
		14'h1e36:	ff_dbi <= 8'h00;
		14'h1e37:	ff_dbi <= 8'h00;
		14'h1e38:	ff_dbi <= 8'h00;
		14'h1e39:	ff_dbi <= 8'h00;
		14'h1e3a:	ff_dbi <= 8'h00;
		14'h1e3b:	ff_dbi <= 8'h00;
		14'h1e3c:	ff_dbi <= 8'h00;
		14'h1e3d:	ff_dbi <= 8'h00;
		14'h1e3e:	ff_dbi <= 8'h00;
		14'h1e3f:	ff_dbi <= 8'h00;
		14'h1e40:	ff_dbi <= 8'h00;
		14'h1e41:	ff_dbi <= 8'h00;
		14'h1e42:	ff_dbi <= 8'h00;
		14'h1e43:	ff_dbi <= 8'h00;
		14'h1e44:	ff_dbi <= 8'h00;
		14'h1e45:	ff_dbi <= 8'h00;
		14'h1e46:	ff_dbi <= 8'h00;
		14'h1e47:	ff_dbi <= 8'h00;
		14'h1e48:	ff_dbi <= 8'h00;
		14'h1e49:	ff_dbi <= 8'h00;
		14'h1e4a:	ff_dbi <= 8'h00;
		14'h1e4b:	ff_dbi <= 8'h00;
		14'h1e4c:	ff_dbi <= 8'h00;
		14'h1e4d:	ff_dbi <= 8'h00;
		14'h1e4e:	ff_dbi <= 8'h00;
		14'h1e4f:	ff_dbi <= 8'h00;
		14'h1e50:	ff_dbi <= 8'h00;
		14'h1e51:	ff_dbi <= 8'h00;
		14'h1e52:	ff_dbi <= 8'h00;
		14'h1e53:	ff_dbi <= 8'h00;
		14'h1e54:	ff_dbi <= 8'h00;
		14'h1e55:	ff_dbi <= 8'h00;
		14'h1e56:	ff_dbi <= 8'h00;
		14'h1e57:	ff_dbi <= 8'h00;
		14'h1e58:	ff_dbi <= 8'h00;
		14'h1e59:	ff_dbi <= 8'h00;
		14'h1e5a:	ff_dbi <= 8'h00;
		14'h1e5b:	ff_dbi <= 8'h00;
		14'h1e5c:	ff_dbi <= 8'h00;
		14'h1e5d:	ff_dbi <= 8'h00;
		14'h1e5e:	ff_dbi <= 8'h00;
		14'h1e5f:	ff_dbi <= 8'h00;
		14'h1e60:	ff_dbi <= 8'h00;
		14'h1e61:	ff_dbi <= 8'h00;
		14'h1e62:	ff_dbi <= 8'h00;
		14'h1e63:	ff_dbi <= 8'h00;
		14'h1e64:	ff_dbi <= 8'h00;
		14'h1e65:	ff_dbi <= 8'h00;
		14'h1e66:	ff_dbi <= 8'h00;
		14'h1e67:	ff_dbi <= 8'h00;
		14'h1e68:	ff_dbi <= 8'h00;
		14'h1e69:	ff_dbi <= 8'h00;
		14'h1e6a:	ff_dbi <= 8'h00;
		14'h1e6b:	ff_dbi <= 8'h00;
		14'h1e6c:	ff_dbi <= 8'h00;
		14'h1e6d:	ff_dbi <= 8'h00;
		14'h1e6e:	ff_dbi <= 8'h00;
		14'h1e6f:	ff_dbi <= 8'h00;
		14'h1e70:	ff_dbi <= 8'h00;
		14'h1e71:	ff_dbi <= 8'h00;
		14'h1e72:	ff_dbi <= 8'h00;
		14'h1e73:	ff_dbi <= 8'h00;
		14'h1e74:	ff_dbi <= 8'h00;
		14'h1e75:	ff_dbi <= 8'h00;
		14'h1e76:	ff_dbi <= 8'h00;
		14'h1e77:	ff_dbi <= 8'h00;
		14'h1e78:	ff_dbi <= 8'h00;
		14'h1e79:	ff_dbi <= 8'h00;
		14'h1e7a:	ff_dbi <= 8'h00;
		14'h1e7b:	ff_dbi <= 8'h00;
		14'h1e7c:	ff_dbi <= 8'h00;
		14'h1e7d:	ff_dbi <= 8'h00;
		14'h1e7e:	ff_dbi <= 8'h00;
		14'h1e7f:	ff_dbi <= 8'h00;
		14'h1e80:	ff_dbi <= 8'h00;
		14'h1e81:	ff_dbi <= 8'h00;
		14'h1e82:	ff_dbi <= 8'h00;
		14'h1e83:	ff_dbi <= 8'h00;
		14'h1e84:	ff_dbi <= 8'h00;
		14'h1e85:	ff_dbi <= 8'h00;
		14'h1e86:	ff_dbi <= 8'h00;
		14'h1e87:	ff_dbi <= 8'h00;
		14'h1e88:	ff_dbi <= 8'h00;
		14'h1e89:	ff_dbi <= 8'h00;
		14'h1e8a:	ff_dbi <= 8'h00;
		14'h1e8b:	ff_dbi <= 8'h00;
		14'h1e8c:	ff_dbi <= 8'h00;
		14'h1e8d:	ff_dbi <= 8'h00;
		14'h1e8e:	ff_dbi <= 8'h00;
		14'h1e8f:	ff_dbi <= 8'h00;
		14'h1e90:	ff_dbi <= 8'h00;
		14'h1e91:	ff_dbi <= 8'h00;
		14'h1e92:	ff_dbi <= 8'h00;
		14'h1e93:	ff_dbi <= 8'h00;
		14'h1e94:	ff_dbi <= 8'h00;
		14'h1e95:	ff_dbi <= 8'h00;
		14'h1e96:	ff_dbi <= 8'h00;
		14'h1e97:	ff_dbi <= 8'h00;
		14'h1e98:	ff_dbi <= 8'h00;
		14'h1e99:	ff_dbi <= 8'h00;
		14'h1e9a:	ff_dbi <= 8'h00;
		14'h1e9b:	ff_dbi <= 8'h00;
		14'h1e9c:	ff_dbi <= 8'h00;
		14'h1e9d:	ff_dbi <= 8'h00;
		14'h1e9e:	ff_dbi <= 8'h00;
		14'h1e9f:	ff_dbi <= 8'h00;
		14'h1ea0:	ff_dbi <= 8'h00;
		14'h1ea1:	ff_dbi <= 8'h00;
		14'h1ea2:	ff_dbi <= 8'h00;
		14'h1ea3:	ff_dbi <= 8'h00;
		14'h1ea4:	ff_dbi <= 8'h00;
		14'h1ea5:	ff_dbi <= 8'h00;
		14'h1ea6:	ff_dbi <= 8'h00;
		14'h1ea7:	ff_dbi <= 8'h00;
		14'h1ea8:	ff_dbi <= 8'h00;
		14'h1ea9:	ff_dbi <= 8'h00;
		14'h1eaa:	ff_dbi <= 8'h00;
		14'h1eab:	ff_dbi <= 8'h00;
		14'h1eac:	ff_dbi <= 8'h00;
		14'h1ead:	ff_dbi <= 8'h00;
		14'h1eae:	ff_dbi <= 8'h00;
		14'h1eaf:	ff_dbi <= 8'h00;
		14'h1eb0:	ff_dbi <= 8'h00;
		14'h1eb1:	ff_dbi <= 8'h00;
		14'h1eb2:	ff_dbi <= 8'h00;
		14'h1eb3:	ff_dbi <= 8'h00;
		14'h1eb4:	ff_dbi <= 8'h00;
		14'h1eb5:	ff_dbi <= 8'h00;
		14'h1eb6:	ff_dbi <= 8'h00;
		14'h1eb7:	ff_dbi <= 8'h00;
		14'h1eb8:	ff_dbi <= 8'h00;
		14'h1eb9:	ff_dbi <= 8'h00;
		14'h1eba:	ff_dbi <= 8'h00;
		14'h1ebb:	ff_dbi <= 8'h00;
		14'h1ebc:	ff_dbi <= 8'h00;
		14'h1ebd:	ff_dbi <= 8'h00;
		14'h1ebe:	ff_dbi <= 8'h00;
		14'h1ebf:	ff_dbi <= 8'h00;
		14'h1ec0:	ff_dbi <= 8'h00;
		14'h1ec1:	ff_dbi <= 8'h00;
		14'h1ec2:	ff_dbi <= 8'h00;
		14'h1ec3:	ff_dbi <= 8'h00;
		14'h1ec4:	ff_dbi <= 8'h00;
		14'h1ec5:	ff_dbi <= 8'h00;
		14'h1ec6:	ff_dbi <= 8'h00;
		14'h1ec7:	ff_dbi <= 8'h00;
		14'h1ec8:	ff_dbi <= 8'h00;
		14'h1ec9:	ff_dbi <= 8'h00;
		14'h1eca:	ff_dbi <= 8'h00;
		14'h1ecb:	ff_dbi <= 8'h00;
		14'h1ecc:	ff_dbi <= 8'h00;
		14'h1ecd:	ff_dbi <= 8'h00;
		14'h1ece:	ff_dbi <= 8'h00;
		14'h1ecf:	ff_dbi <= 8'h00;
		14'h1ed0:	ff_dbi <= 8'h00;
		14'h1ed1:	ff_dbi <= 8'h00;
		14'h1ed2:	ff_dbi <= 8'h00;
		14'h1ed3:	ff_dbi <= 8'h00;
		14'h1ed4:	ff_dbi <= 8'h00;
		14'h1ed5:	ff_dbi <= 8'h00;
		14'h1ed6:	ff_dbi <= 8'h00;
		14'h1ed7:	ff_dbi <= 8'h00;
		14'h1ed8:	ff_dbi <= 8'h00;
		14'h1ed9:	ff_dbi <= 8'h00;
		14'h1eda:	ff_dbi <= 8'h00;
		14'h1edb:	ff_dbi <= 8'h00;
		14'h1edc:	ff_dbi <= 8'h00;
		14'h1edd:	ff_dbi <= 8'h00;
		14'h1ede:	ff_dbi <= 8'h00;
		14'h1edf:	ff_dbi <= 8'h00;
		14'h1ee0:	ff_dbi <= 8'h00;
		14'h1ee1:	ff_dbi <= 8'h00;
		14'h1ee2:	ff_dbi <= 8'h00;
		14'h1ee3:	ff_dbi <= 8'h00;
		14'h1ee4:	ff_dbi <= 8'h00;
		14'h1ee5:	ff_dbi <= 8'h00;
		14'h1ee6:	ff_dbi <= 8'h00;
		14'h1ee7:	ff_dbi <= 8'h00;
		14'h1ee8:	ff_dbi <= 8'h00;
		14'h1ee9:	ff_dbi <= 8'h00;
		14'h1eea:	ff_dbi <= 8'h00;
		14'h1eeb:	ff_dbi <= 8'h00;
		14'h1eec:	ff_dbi <= 8'h00;
		14'h1eed:	ff_dbi <= 8'h00;
		14'h1eee:	ff_dbi <= 8'h00;
		14'h1eef:	ff_dbi <= 8'h00;
		14'h1ef0:	ff_dbi <= 8'h00;
		14'h1ef1:	ff_dbi <= 8'h00;
		14'h1ef2:	ff_dbi <= 8'h00;
		14'h1ef3:	ff_dbi <= 8'h00;
		14'h1ef4:	ff_dbi <= 8'h00;
		14'h1ef5:	ff_dbi <= 8'h00;
		14'h1ef6:	ff_dbi <= 8'h00;
		14'h1ef7:	ff_dbi <= 8'h00;
		14'h1ef8:	ff_dbi <= 8'h00;
		14'h1ef9:	ff_dbi <= 8'h00;
		14'h1efa:	ff_dbi <= 8'h00;
		14'h1efb:	ff_dbi <= 8'h00;
		14'h1efc:	ff_dbi <= 8'h00;
		14'h1efd:	ff_dbi <= 8'h00;
		14'h1efe:	ff_dbi <= 8'h00;
		14'h1eff:	ff_dbi <= 8'h00;
		14'h1f00:	ff_dbi <= 8'h00;
		14'h1f01:	ff_dbi <= 8'h00;
		14'h1f02:	ff_dbi <= 8'h00;
		14'h1f03:	ff_dbi <= 8'h00;
		14'h1f04:	ff_dbi <= 8'h00;
		14'h1f05:	ff_dbi <= 8'h00;
		14'h1f06:	ff_dbi <= 8'h00;
		14'h1f07:	ff_dbi <= 8'h00;
		14'h1f08:	ff_dbi <= 8'h00;
		14'h1f09:	ff_dbi <= 8'h00;
		14'h1f0a:	ff_dbi <= 8'h00;
		14'h1f0b:	ff_dbi <= 8'h00;
		14'h1f0c:	ff_dbi <= 8'h00;
		14'h1f0d:	ff_dbi <= 8'h00;
		14'h1f0e:	ff_dbi <= 8'h00;
		14'h1f0f:	ff_dbi <= 8'h00;
		14'h1f10:	ff_dbi <= 8'h00;
		14'h1f11:	ff_dbi <= 8'h00;
		14'h1f12:	ff_dbi <= 8'h00;
		14'h1f13:	ff_dbi <= 8'h00;
		14'h1f14:	ff_dbi <= 8'h00;
		14'h1f15:	ff_dbi <= 8'h00;
		14'h1f16:	ff_dbi <= 8'h00;
		14'h1f17:	ff_dbi <= 8'h00;
		14'h1f18:	ff_dbi <= 8'h00;
		14'h1f19:	ff_dbi <= 8'h00;
		14'h1f1a:	ff_dbi <= 8'h00;
		14'h1f1b:	ff_dbi <= 8'h00;
		14'h1f1c:	ff_dbi <= 8'h00;
		14'h1f1d:	ff_dbi <= 8'h00;
		14'h1f1e:	ff_dbi <= 8'h00;
		14'h1f1f:	ff_dbi <= 8'h00;
		14'h1f20:	ff_dbi <= 8'h00;
		14'h1f21:	ff_dbi <= 8'h00;
		14'h1f22:	ff_dbi <= 8'h00;
		14'h1f23:	ff_dbi <= 8'h00;
		14'h1f24:	ff_dbi <= 8'h00;
		14'h1f25:	ff_dbi <= 8'h00;
		14'h1f26:	ff_dbi <= 8'h00;
		14'h1f27:	ff_dbi <= 8'h00;
		14'h1f28:	ff_dbi <= 8'h00;
		14'h1f29:	ff_dbi <= 8'h00;
		14'h1f2a:	ff_dbi <= 8'h00;
		14'h1f2b:	ff_dbi <= 8'h00;
		14'h1f2c:	ff_dbi <= 8'h00;
		14'h1f2d:	ff_dbi <= 8'h00;
		14'h1f2e:	ff_dbi <= 8'h00;
		14'h1f2f:	ff_dbi <= 8'h00;
		14'h1f30:	ff_dbi <= 8'h00;
		14'h1f31:	ff_dbi <= 8'h00;
		14'h1f32:	ff_dbi <= 8'h00;
		14'h1f33:	ff_dbi <= 8'h00;
		14'h1f34:	ff_dbi <= 8'h00;
		14'h1f35:	ff_dbi <= 8'h00;
		14'h1f36:	ff_dbi <= 8'h00;
		14'h1f37:	ff_dbi <= 8'h00;
		14'h1f38:	ff_dbi <= 8'h00;
		14'h1f39:	ff_dbi <= 8'h00;
		14'h1f3a:	ff_dbi <= 8'h00;
		14'h1f3b:	ff_dbi <= 8'h00;
		14'h1f3c:	ff_dbi <= 8'h00;
		14'h1f3d:	ff_dbi <= 8'h00;
		14'h1f3e:	ff_dbi <= 8'h00;
		14'h1f3f:	ff_dbi <= 8'h00;
		14'h1f40:	ff_dbi <= 8'h00;
		14'h1f41:	ff_dbi <= 8'h00;
		14'h1f42:	ff_dbi <= 8'h00;
		14'h1f43:	ff_dbi <= 8'h00;
		14'h1f44:	ff_dbi <= 8'h00;
		14'h1f45:	ff_dbi <= 8'h00;
		14'h1f46:	ff_dbi <= 8'h00;
		14'h1f47:	ff_dbi <= 8'h00;
		14'h1f48:	ff_dbi <= 8'h00;
		14'h1f49:	ff_dbi <= 8'h00;
		14'h1f4a:	ff_dbi <= 8'h00;
		14'h1f4b:	ff_dbi <= 8'h00;
		14'h1f4c:	ff_dbi <= 8'h00;
		14'h1f4d:	ff_dbi <= 8'h00;
		14'h1f4e:	ff_dbi <= 8'h00;
		14'h1f4f:	ff_dbi <= 8'h00;
		14'h1f50:	ff_dbi <= 8'h00;
		14'h1f51:	ff_dbi <= 8'h00;
		14'h1f52:	ff_dbi <= 8'h00;
		14'h1f53:	ff_dbi <= 8'h00;
		14'h1f54:	ff_dbi <= 8'h00;
		14'h1f55:	ff_dbi <= 8'h00;
		14'h1f56:	ff_dbi <= 8'h00;
		14'h1f57:	ff_dbi <= 8'h00;
		14'h1f58:	ff_dbi <= 8'h00;
		14'h1f59:	ff_dbi <= 8'h00;
		14'h1f5a:	ff_dbi <= 8'h00;
		14'h1f5b:	ff_dbi <= 8'h00;
		14'h1f5c:	ff_dbi <= 8'h00;
		14'h1f5d:	ff_dbi <= 8'h00;
		14'h1f5e:	ff_dbi <= 8'h00;
		14'h1f5f:	ff_dbi <= 8'h00;
		14'h1f60:	ff_dbi <= 8'h00;
		14'h1f61:	ff_dbi <= 8'h00;
		14'h1f62:	ff_dbi <= 8'h00;
		14'h1f63:	ff_dbi <= 8'h00;
		14'h1f64:	ff_dbi <= 8'h00;
		14'h1f65:	ff_dbi <= 8'h00;
		14'h1f66:	ff_dbi <= 8'h00;
		14'h1f67:	ff_dbi <= 8'h00;
		14'h1f68:	ff_dbi <= 8'h00;
		14'h1f69:	ff_dbi <= 8'h00;
		14'h1f6a:	ff_dbi <= 8'h00;
		14'h1f6b:	ff_dbi <= 8'h00;
		14'h1f6c:	ff_dbi <= 8'h00;
		14'h1f6d:	ff_dbi <= 8'h00;
		14'h1f6e:	ff_dbi <= 8'h00;
		14'h1f6f:	ff_dbi <= 8'h00;
		14'h1f70:	ff_dbi <= 8'h00;
		14'h1f71:	ff_dbi <= 8'h00;
		14'h1f72:	ff_dbi <= 8'h00;
		14'h1f73:	ff_dbi <= 8'h00;
		14'h1f74:	ff_dbi <= 8'h00;
		14'h1f75:	ff_dbi <= 8'h00;
		14'h1f76:	ff_dbi <= 8'h00;
		14'h1f77:	ff_dbi <= 8'h00;
		14'h1f78:	ff_dbi <= 8'h00;
		14'h1f79:	ff_dbi <= 8'h00;
		14'h1f7a:	ff_dbi <= 8'h00;
		14'h1f7b:	ff_dbi <= 8'h00;
		14'h1f7c:	ff_dbi <= 8'h00;
		14'h1f7d:	ff_dbi <= 8'h00;
		14'h1f7e:	ff_dbi <= 8'h00;
		14'h1f7f:	ff_dbi <= 8'h00;
		14'h1f80:	ff_dbi <= 8'h00;
		14'h1f81:	ff_dbi <= 8'h00;
		14'h1f82:	ff_dbi <= 8'h00;
		14'h1f83:	ff_dbi <= 8'h00;
		14'h1f84:	ff_dbi <= 8'h00;
		14'h1f85:	ff_dbi <= 8'h00;
		14'h1f86:	ff_dbi <= 8'h00;
		14'h1f87:	ff_dbi <= 8'h00;
		14'h1f88:	ff_dbi <= 8'h00;
		14'h1f89:	ff_dbi <= 8'h00;
		14'h1f8a:	ff_dbi <= 8'h00;
		14'h1f8b:	ff_dbi <= 8'h00;
		14'h1f8c:	ff_dbi <= 8'h00;
		14'h1f8d:	ff_dbi <= 8'h00;
		14'h1f8e:	ff_dbi <= 8'h00;
		14'h1f8f:	ff_dbi <= 8'h00;
		14'h1f90:	ff_dbi <= 8'h00;
		14'h1f91:	ff_dbi <= 8'h00;
		14'h1f92:	ff_dbi <= 8'h00;
		14'h1f93:	ff_dbi <= 8'h00;
		14'h1f94:	ff_dbi <= 8'h00;
		14'h1f95:	ff_dbi <= 8'h00;
		14'h1f96:	ff_dbi <= 8'h00;
		14'h1f97:	ff_dbi <= 8'h00;
		14'h1f98:	ff_dbi <= 8'h00;
		14'h1f99:	ff_dbi <= 8'h00;
		14'h1f9a:	ff_dbi <= 8'h00;
		14'h1f9b:	ff_dbi <= 8'h00;
		14'h1f9c:	ff_dbi <= 8'h00;
		14'h1f9d:	ff_dbi <= 8'h00;
		14'h1f9e:	ff_dbi <= 8'h00;
		14'h1f9f:	ff_dbi <= 8'h00;
		14'h1fa0:	ff_dbi <= 8'h00;
		14'h1fa1:	ff_dbi <= 8'h00;
		14'h1fa2:	ff_dbi <= 8'h00;
		14'h1fa3:	ff_dbi <= 8'h00;
		14'h1fa4:	ff_dbi <= 8'h00;
		14'h1fa5:	ff_dbi <= 8'h00;
		14'h1fa6:	ff_dbi <= 8'h00;
		14'h1fa7:	ff_dbi <= 8'h00;
		14'h1fa8:	ff_dbi <= 8'h00;
		14'h1fa9:	ff_dbi <= 8'h00;
		14'h1faa:	ff_dbi <= 8'h00;
		14'h1fab:	ff_dbi <= 8'h00;
		14'h1fac:	ff_dbi <= 8'h00;
		14'h1fad:	ff_dbi <= 8'h00;
		14'h1fae:	ff_dbi <= 8'h00;
		14'h1faf:	ff_dbi <= 8'h00;
		14'h1fb0:	ff_dbi <= 8'h00;
		14'h1fb1:	ff_dbi <= 8'h00;
		14'h1fb2:	ff_dbi <= 8'h00;
		14'h1fb3:	ff_dbi <= 8'h00;
		14'h1fb4:	ff_dbi <= 8'h00;
		14'h1fb5:	ff_dbi <= 8'h00;
		14'h1fb6:	ff_dbi <= 8'h00;
		14'h1fb7:	ff_dbi <= 8'h00;
		14'h1fb8:	ff_dbi <= 8'h00;
		14'h1fb9:	ff_dbi <= 8'h00;
		14'h1fba:	ff_dbi <= 8'h00;
		14'h1fbb:	ff_dbi <= 8'h00;
		14'h1fbc:	ff_dbi <= 8'h00;
		14'h1fbd:	ff_dbi <= 8'h00;
		14'h1fbe:	ff_dbi <= 8'h00;
		14'h1fbf:	ff_dbi <= 8'h00;
		14'h1fc0:	ff_dbi <= 8'h00;
		14'h1fc1:	ff_dbi <= 8'h00;
		14'h1fc2:	ff_dbi <= 8'h00;
		14'h1fc3:	ff_dbi <= 8'h00;
		14'h1fc4:	ff_dbi <= 8'h00;
		14'h1fc5:	ff_dbi <= 8'h00;
		14'h1fc6:	ff_dbi <= 8'h00;
		14'h1fc7:	ff_dbi <= 8'h00;
		14'h1fc8:	ff_dbi <= 8'h00;
		14'h1fc9:	ff_dbi <= 8'h00;
		14'h1fca:	ff_dbi <= 8'h00;
		14'h1fcb:	ff_dbi <= 8'h00;
		14'h1fcc:	ff_dbi <= 8'h00;
		14'h1fcd:	ff_dbi <= 8'h00;
		14'h1fce:	ff_dbi <= 8'h00;
		14'h1fcf:	ff_dbi <= 8'h00;
		14'h1fd0:	ff_dbi <= 8'h00;
		14'h1fd1:	ff_dbi <= 8'h00;
		14'h1fd2:	ff_dbi <= 8'h00;
		14'h1fd3:	ff_dbi <= 8'h00;
		14'h1fd4:	ff_dbi <= 8'h00;
		14'h1fd5:	ff_dbi <= 8'h00;
		14'h1fd6:	ff_dbi <= 8'h00;
		14'h1fd7:	ff_dbi <= 8'h00;
		14'h1fd8:	ff_dbi <= 8'h00;
		14'h1fd9:	ff_dbi <= 8'h00;
		14'h1fda:	ff_dbi <= 8'h00;
		14'h1fdb:	ff_dbi <= 8'h00;
		14'h1fdc:	ff_dbi <= 8'h00;
		14'h1fdd:	ff_dbi <= 8'h00;
		14'h1fde:	ff_dbi <= 8'h00;
		14'h1fdf:	ff_dbi <= 8'h00;
		14'h1fe0:	ff_dbi <= 8'h00;
		14'h1fe1:	ff_dbi <= 8'h00;
		14'h1fe2:	ff_dbi <= 8'h00;
		14'h1fe3:	ff_dbi <= 8'h00;
		14'h1fe4:	ff_dbi <= 8'h00;
		14'h1fe5:	ff_dbi <= 8'h00;
		14'h1fe6:	ff_dbi <= 8'h00;
		14'h1fe7:	ff_dbi <= 8'h00;
		14'h1fe8:	ff_dbi <= 8'h00;
		14'h1fe9:	ff_dbi <= 8'h00;
		14'h1fea:	ff_dbi <= 8'h00;
		14'h1feb:	ff_dbi <= 8'h00;
		14'h1fec:	ff_dbi <= 8'h00;
		14'h1fed:	ff_dbi <= 8'h00;
		14'h1fee:	ff_dbi <= 8'h00;
		14'h1fef:	ff_dbi <= 8'h00;
		14'h1ff0:	ff_dbi <= 8'h00;
		14'h1ff1:	ff_dbi <= 8'h00;
		14'h1ff2:	ff_dbi <= 8'h00;
		14'h1ff3:	ff_dbi <= 8'h00;
		14'h1ff4:	ff_dbi <= 8'h00;
		14'h1ff5:	ff_dbi <= 8'h00;
		14'h1ff6:	ff_dbi <= 8'h00;
		14'h1ff7:	ff_dbi <= 8'h00;
		14'h1ff8:	ff_dbi <= 8'h00;
		14'h1ff9:	ff_dbi <= 8'h00;
		14'h1ffa:	ff_dbi <= 8'h00;
		14'h1ffb:	ff_dbi <= 8'h00;
		14'h1ffc:	ff_dbi <= 8'h00;
		14'h1ffd:	ff_dbi <= 8'h00;
		14'h1ffe:	ff_dbi <= 8'h00;
		14'h1fff:	ff_dbi <= 8'h00;
		14'h2000:	ff_dbi <= 8'hf4;
		14'h2001:	ff_dbi <= 8'hf4;
		14'h2002:	ff_dbi <= 8'hf4;
		14'h2003:	ff_dbi <= 8'hf4;
		14'h2004:	ff_dbi <= 8'hf4;
		14'h2005:	ff_dbi <= 8'hf4;
		14'h2006:	ff_dbi <= 8'hf4;
		14'h2007:	ff_dbi <= 8'hf4;
		14'h2008:	ff_dbi <= 8'hf4;
		14'h2009:	ff_dbi <= 8'hf4;
		14'h200a:	ff_dbi <= 8'hf4;
		14'h200b:	ff_dbi <= 8'hf4;
		14'h200c:	ff_dbi <= 8'hf4;
		14'h200d:	ff_dbi <= 8'hf4;
		14'h200e:	ff_dbi <= 8'hf4;
		14'h200f:	ff_dbi <= 8'hf4;
		14'h2010:	ff_dbi <= 8'hf4;
		14'h2011:	ff_dbi <= 8'hf4;
		14'h2012:	ff_dbi <= 8'hf4;
		14'h2013:	ff_dbi <= 8'hf4;
		14'h2014:	ff_dbi <= 8'hf4;
		14'h2015:	ff_dbi <= 8'hf4;
		14'h2016:	ff_dbi <= 8'hf4;
		14'h2017:	ff_dbi <= 8'hf4;
		14'h2018:	ff_dbi <= 8'hf4;
		14'h2019:	ff_dbi <= 8'hf4;
		14'h201a:	ff_dbi <= 8'hf4;
		14'h201b:	ff_dbi <= 8'hf4;
		14'h201c:	ff_dbi <= 8'hf4;
		14'h201d:	ff_dbi <= 8'hf4;
		14'h201e:	ff_dbi <= 8'hf4;
		14'h201f:	ff_dbi <= 8'hf4;
		14'h2020:	ff_dbi <= 8'h00;
		14'h2021:	ff_dbi <= 8'h00;
		14'h2022:	ff_dbi <= 8'h00;
		14'h2023:	ff_dbi <= 8'h00;
		14'h2024:	ff_dbi <= 8'h11;
		14'h2025:	ff_dbi <= 8'h06;
		14'h2026:	ff_dbi <= 8'h33;
		14'h2027:	ff_dbi <= 8'h07;
		14'h2028:	ff_dbi <= 8'h17;
		14'h2029:	ff_dbi <= 8'h01;
		14'h202a:	ff_dbi <= 8'h27;
		14'h202b:	ff_dbi <= 8'h03;
		14'h202c:	ff_dbi <= 8'h51;
		14'h202d:	ff_dbi <= 8'h01;
		14'h202e:	ff_dbi <= 8'h27;
		14'h202f:	ff_dbi <= 8'h06;
		14'h2030:	ff_dbi <= 8'h71;
		14'h2031:	ff_dbi <= 8'h01;
		14'h2032:	ff_dbi <= 8'h73;
		14'h2033:	ff_dbi <= 8'h03;
		14'h2034:	ff_dbi <= 8'h61;
		14'h2035:	ff_dbi <= 8'h06;
		14'h2036:	ff_dbi <= 8'h64;
		14'h2037:	ff_dbi <= 8'h06;
		14'h2038:	ff_dbi <= 8'h11;
		14'h2039:	ff_dbi <= 8'h04;
		14'h203a:	ff_dbi <= 8'h65;
		14'h203b:	ff_dbi <= 8'h02;
		14'h203c:	ff_dbi <= 8'h55;
		14'h203d:	ff_dbi <= 8'h05;
		14'h203e:	ff_dbi <= 8'h77;
		14'h203f:	ff_dbi <= 8'h07;
		14'h2040:	ff_dbi <= 8'h00;
		14'h2041:	ff_dbi <= 8'h00;
		14'h2042:	ff_dbi <= 8'h00;
		14'h2043:	ff_dbi <= 8'h00;
		14'h2044:	ff_dbi <= 8'h00;
		14'h2045:	ff_dbi <= 8'h00;
		14'h2046:	ff_dbi <= 8'h00;
		14'h2047:	ff_dbi <= 8'h00;
		14'h2048:	ff_dbi <= 8'h00;
		14'h2049:	ff_dbi <= 8'h00;
		14'h204a:	ff_dbi <= 8'h00;
		14'h204b:	ff_dbi <= 8'h00;
		14'h204c:	ff_dbi <= 8'h00;
		14'h204d:	ff_dbi <= 8'h00;
		14'h204e:	ff_dbi <= 8'h00;
		14'h204f:	ff_dbi <= 8'h00;
		14'h2050:	ff_dbi <= 8'h00;
		14'h2051:	ff_dbi <= 8'h00;
		14'h2052:	ff_dbi <= 8'h00;
		14'h2053:	ff_dbi <= 8'h00;
		14'h2054:	ff_dbi <= 8'h00;
		14'h2055:	ff_dbi <= 8'h00;
		14'h2056:	ff_dbi <= 8'h00;
		14'h2057:	ff_dbi <= 8'h00;
		14'h2058:	ff_dbi <= 8'h00;
		14'h2059:	ff_dbi <= 8'h00;
		14'h205a:	ff_dbi <= 8'h00;
		14'h205b:	ff_dbi <= 8'h00;
		14'h205c:	ff_dbi <= 8'h00;
		14'h205d:	ff_dbi <= 8'h00;
		14'h205e:	ff_dbi <= 8'h00;
		14'h205f:	ff_dbi <= 8'h00;
		14'h2060:	ff_dbi <= 8'h00;
		14'h2061:	ff_dbi <= 8'h00;
		14'h2062:	ff_dbi <= 8'h00;
		14'h2063:	ff_dbi <= 8'h00;
		14'h2064:	ff_dbi <= 8'h00;
		14'h2065:	ff_dbi <= 8'h00;
		14'h2066:	ff_dbi <= 8'h00;
		14'h2067:	ff_dbi <= 8'h00;
		14'h2068:	ff_dbi <= 8'h00;
		14'h2069:	ff_dbi <= 8'h00;
		14'h206a:	ff_dbi <= 8'h00;
		14'h206b:	ff_dbi <= 8'h00;
		14'h206c:	ff_dbi <= 8'h00;
		14'h206d:	ff_dbi <= 8'h00;
		14'h206e:	ff_dbi <= 8'h00;
		14'h206f:	ff_dbi <= 8'h00;
		14'h2070:	ff_dbi <= 8'h00;
		14'h2071:	ff_dbi <= 8'h00;
		14'h2072:	ff_dbi <= 8'h00;
		14'h2073:	ff_dbi <= 8'h00;
		14'h2074:	ff_dbi <= 8'h00;
		14'h2075:	ff_dbi <= 8'h00;
		14'h2076:	ff_dbi <= 8'h00;
		14'h2077:	ff_dbi <= 8'h00;
		14'h2078:	ff_dbi <= 8'h00;
		14'h2079:	ff_dbi <= 8'h00;
		14'h207a:	ff_dbi <= 8'h00;
		14'h207b:	ff_dbi <= 8'h00;
		14'h207c:	ff_dbi <= 8'h00;
		14'h207d:	ff_dbi <= 8'h00;
		14'h207e:	ff_dbi <= 8'h00;
		14'h207f:	ff_dbi <= 8'h00;
		14'h2080:	ff_dbi <= 8'h00;
		14'h2081:	ff_dbi <= 8'h00;
		14'h2082:	ff_dbi <= 8'h00;
		14'h2083:	ff_dbi <= 8'h00;
		14'h2084:	ff_dbi <= 8'h00;
		14'h2085:	ff_dbi <= 8'h00;
		14'h2086:	ff_dbi <= 8'h00;
		14'h2087:	ff_dbi <= 8'h00;
		14'h2088:	ff_dbi <= 8'h00;
		14'h2089:	ff_dbi <= 8'h00;
		14'h208a:	ff_dbi <= 8'h00;
		14'h208b:	ff_dbi <= 8'h00;
		14'h208c:	ff_dbi <= 8'h00;
		14'h208d:	ff_dbi <= 8'h00;
		14'h208e:	ff_dbi <= 8'h00;
		14'h208f:	ff_dbi <= 8'h00;
		14'h2090:	ff_dbi <= 8'h00;
		14'h2091:	ff_dbi <= 8'h00;
		14'h2092:	ff_dbi <= 8'h00;
		14'h2093:	ff_dbi <= 8'h00;
		14'h2094:	ff_dbi <= 8'h00;
		14'h2095:	ff_dbi <= 8'h00;
		14'h2096:	ff_dbi <= 8'h00;
		14'h2097:	ff_dbi <= 8'h00;
		14'h2098:	ff_dbi <= 8'h00;
		14'h2099:	ff_dbi <= 8'h00;
		14'h209a:	ff_dbi <= 8'h00;
		14'h209b:	ff_dbi <= 8'h00;
		14'h209c:	ff_dbi <= 8'h00;
		14'h209d:	ff_dbi <= 8'h00;
		14'h209e:	ff_dbi <= 8'h00;
		14'h209f:	ff_dbi <= 8'h00;
		14'h20a0:	ff_dbi <= 8'h00;
		14'h20a1:	ff_dbi <= 8'h00;
		14'h20a2:	ff_dbi <= 8'h00;
		14'h20a3:	ff_dbi <= 8'h00;
		14'h20a4:	ff_dbi <= 8'h00;
		14'h20a5:	ff_dbi <= 8'h00;
		14'h20a6:	ff_dbi <= 8'h00;
		14'h20a7:	ff_dbi <= 8'h00;
		14'h20a8:	ff_dbi <= 8'h00;
		14'h20a9:	ff_dbi <= 8'h00;
		14'h20aa:	ff_dbi <= 8'h00;
		14'h20ab:	ff_dbi <= 8'h00;
		14'h20ac:	ff_dbi <= 8'h00;
		14'h20ad:	ff_dbi <= 8'h00;
		14'h20ae:	ff_dbi <= 8'h00;
		14'h20af:	ff_dbi <= 8'h00;
		14'h20b0:	ff_dbi <= 8'h00;
		14'h20b1:	ff_dbi <= 8'h00;
		14'h20b2:	ff_dbi <= 8'h00;
		14'h20b3:	ff_dbi <= 8'h00;
		14'h20b4:	ff_dbi <= 8'h00;
		14'h20b5:	ff_dbi <= 8'h00;
		14'h20b6:	ff_dbi <= 8'h00;
		14'h20b7:	ff_dbi <= 8'h00;
		14'h20b8:	ff_dbi <= 8'h00;
		14'h20b9:	ff_dbi <= 8'h00;
		14'h20ba:	ff_dbi <= 8'h00;
		14'h20bb:	ff_dbi <= 8'h00;
		14'h20bc:	ff_dbi <= 8'h00;
		14'h20bd:	ff_dbi <= 8'h00;
		14'h20be:	ff_dbi <= 8'h00;
		14'h20bf:	ff_dbi <= 8'h00;
		14'h20c0:	ff_dbi <= 8'h00;
		14'h20c1:	ff_dbi <= 8'h00;
		14'h20c2:	ff_dbi <= 8'h00;
		14'h20c3:	ff_dbi <= 8'h00;
		14'h20c4:	ff_dbi <= 8'h00;
		14'h20c5:	ff_dbi <= 8'h00;
		14'h20c6:	ff_dbi <= 8'h00;
		14'h20c7:	ff_dbi <= 8'h00;
		14'h20c8:	ff_dbi <= 8'h00;
		14'h20c9:	ff_dbi <= 8'h00;
		14'h20ca:	ff_dbi <= 8'h00;
		14'h20cb:	ff_dbi <= 8'h00;
		14'h20cc:	ff_dbi <= 8'h00;
		14'h20cd:	ff_dbi <= 8'h00;
		14'h20ce:	ff_dbi <= 8'h00;
		14'h20cf:	ff_dbi <= 8'h00;
		14'h20d0:	ff_dbi <= 8'h00;
		14'h20d1:	ff_dbi <= 8'h00;
		14'h20d2:	ff_dbi <= 8'h00;
		14'h20d3:	ff_dbi <= 8'h00;
		14'h20d4:	ff_dbi <= 8'h00;
		14'h20d5:	ff_dbi <= 8'h00;
		14'h20d6:	ff_dbi <= 8'h00;
		14'h20d7:	ff_dbi <= 8'h00;
		14'h20d8:	ff_dbi <= 8'h00;
		14'h20d9:	ff_dbi <= 8'h00;
		14'h20da:	ff_dbi <= 8'h00;
		14'h20db:	ff_dbi <= 8'h00;
		14'h20dc:	ff_dbi <= 8'h00;
		14'h20dd:	ff_dbi <= 8'h00;
		14'h20de:	ff_dbi <= 8'h00;
		14'h20df:	ff_dbi <= 8'h00;
		14'h20e0:	ff_dbi <= 8'h00;
		14'h20e1:	ff_dbi <= 8'h00;
		14'h20e2:	ff_dbi <= 8'h00;
		14'h20e3:	ff_dbi <= 8'h00;
		14'h20e4:	ff_dbi <= 8'h00;
		14'h20e5:	ff_dbi <= 8'h00;
		14'h20e6:	ff_dbi <= 8'h00;
		14'h20e7:	ff_dbi <= 8'h00;
		14'h20e8:	ff_dbi <= 8'h00;
		14'h20e9:	ff_dbi <= 8'h00;
		14'h20ea:	ff_dbi <= 8'h00;
		14'h20eb:	ff_dbi <= 8'h00;
		14'h20ec:	ff_dbi <= 8'h00;
		14'h20ed:	ff_dbi <= 8'h00;
		14'h20ee:	ff_dbi <= 8'h00;
		14'h20ef:	ff_dbi <= 8'h00;
		14'h20f0:	ff_dbi <= 8'h00;
		14'h20f1:	ff_dbi <= 8'h00;
		14'h20f2:	ff_dbi <= 8'h00;
		14'h20f3:	ff_dbi <= 8'h00;
		14'h20f4:	ff_dbi <= 8'h00;
		14'h20f5:	ff_dbi <= 8'h00;
		14'h20f6:	ff_dbi <= 8'h00;
		14'h20f7:	ff_dbi <= 8'h00;
		14'h20f8:	ff_dbi <= 8'h00;
		14'h20f9:	ff_dbi <= 8'h00;
		14'h20fa:	ff_dbi <= 8'h00;
		14'h20fb:	ff_dbi <= 8'h00;
		14'h20fc:	ff_dbi <= 8'h00;
		14'h20fd:	ff_dbi <= 8'h00;
		14'h20fe:	ff_dbi <= 8'h00;
		14'h20ff:	ff_dbi <= 8'h00;
		14'h2100:	ff_dbi <= 8'h00;
		14'h2101:	ff_dbi <= 8'h00;
		14'h2102:	ff_dbi <= 8'h00;
		14'h2103:	ff_dbi <= 8'h00;
		14'h2104:	ff_dbi <= 8'h00;
		14'h2105:	ff_dbi <= 8'h00;
		14'h2106:	ff_dbi <= 8'h00;
		14'h2107:	ff_dbi <= 8'h00;
		14'h2108:	ff_dbi <= 8'h00;
		14'h2109:	ff_dbi <= 8'h00;
		14'h210a:	ff_dbi <= 8'h00;
		14'h210b:	ff_dbi <= 8'h00;
		14'h210c:	ff_dbi <= 8'h00;
		14'h210d:	ff_dbi <= 8'h00;
		14'h210e:	ff_dbi <= 8'h00;
		14'h210f:	ff_dbi <= 8'h00;
		14'h2110:	ff_dbi <= 8'h00;
		14'h2111:	ff_dbi <= 8'h00;
		14'h2112:	ff_dbi <= 8'h00;
		14'h2113:	ff_dbi <= 8'h00;
		14'h2114:	ff_dbi <= 8'h00;
		14'h2115:	ff_dbi <= 8'h00;
		14'h2116:	ff_dbi <= 8'h00;
		14'h2117:	ff_dbi <= 8'h00;
		14'h2118:	ff_dbi <= 8'h00;
		14'h2119:	ff_dbi <= 8'h00;
		14'h211a:	ff_dbi <= 8'h00;
		14'h211b:	ff_dbi <= 8'h00;
		14'h211c:	ff_dbi <= 8'h00;
		14'h211d:	ff_dbi <= 8'h00;
		14'h211e:	ff_dbi <= 8'h00;
		14'h211f:	ff_dbi <= 8'h00;
		14'h2120:	ff_dbi <= 8'h00;
		14'h2121:	ff_dbi <= 8'h00;
		14'h2122:	ff_dbi <= 8'h00;
		14'h2123:	ff_dbi <= 8'h00;
		14'h2124:	ff_dbi <= 8'h00;
		14'h2125:	ff_dbi <= 8'h00;
		14'h2126:	ff_dbi <= 8'h00;
		14'h2127:	ff_dbi <= 8'h00;
		14'h2128:	ff_dbi <= 8'h00;
		14'h2129:	ff_dbi <= 8'h00;
		14'h212a:	ff_dbi <= 8'h00;
		14'h212b:	ff_dbi <= 8'h00;
		14'h212c:	ff_dbi <= 8'h00;
		14'h212d:	ff_dbi <= 8'h00;
		14'h212e:	ff_dbi <= 8'h00;
		14'h212f:	ff_dbi <= 8'h00;
		14'h2130:	ff_dbi <= 8'h00;
		14'h2131:	ff_dbi <= 8'h00;
		14'h2132:	ff_dbi <= 8'h00;
		14'h2133:	ff_dbi <= 8'h00;
		14'h2134:	ff_dbi <= 8'h00;
		14'h2135:	ff_dbi <= 8'h00;
		14'h2136:	ff_dbi <= 8'h00;
		14'h2137:	ff_dbi <= 8'h00;
		14'h2138:	ff_dbi <= 8'h00;
		14'h2139:	ff_dbi <= 8'h00;
		14'h213a:	ff_dbi <= 8'h00;
		14'h213b:	ff_dbi <= 8'h00;
		14'h213c:	ff_dbi <= 8'h00;
		14'h213d:	ff_dbi <= 8'h00;
		14'h213e:	ff_dbi <= 8'h00;
		14'h213f:	ff_dbi <= 8'h00;
		14'h2140:	ff_dbi <= 8'h00;
		14'h2141:	ff_dbi <= 8'h00;
		14'h2142:	ff_dbi <= 8'h00;
		14'h2143:	ff_dbi <= 8'h00;
		14'h2144:	ff_dbi <= 8'h00;
		14'h2145:	ff_dbi <= 8'h00;
		14'h2146:	ff_dbi <= 8'h00;
		14'h2147:	ff_dbi <= 8'h00;
		14'h2148:	ff_dbi <= 8'h00;
		14'h2149:	ff_dbi <= 8'h00;
		14'h214a:	ff_dbi <= 8'h00;
		14'h214b:	ff_dbi <= 8'h00;
		14'h214c:	ff_dbi <= 8'h00;
		14'h214d:	ff_dbi <= 8'h00;
		14'h214e:	ff_dbi <= 8'h00;
		14'h214f:	ff_dbi <= 8'h00;
		14'h2150:	ff_dbi <= 8'h00;
		14'h2151:	ff_dbi <= 8'h00;
		14'h2152:	ff_dbi <= 8'h00;
		14'h2153:	ff_dbi <= 8'h00;
		14'h2154:	ff_dbi <= 8'h00;
		14'h2155:	ff_dbi <= 8'h00;
		14'h2156:	ff_dbi <= 8'h00;
		14'h2157:	ff_dbi <= 8'h00;
		14'h2158:	ff_dbi <= 8'h00;
		14'h2159:	ff_dbi <= 8'h00;
		14'h215a:	ff_dbi <= 8'h00;
		14'h215b:	ff_dbi <= 8'h00;
		14'h215c:	ff_dbi <= 8'h00;
		14'h215d:	ff_dbi <= 8'h00;
		14'h215e:	ff_dbi <= 8'h00;
		14'h215f:	ff_dbi <= 8'h00;
		14'h2160:	ff_dbi <= 8'h00;
		14'h2161:	ff_dbi <= 8'h00;
		14'h2162:	ff_dbi <= 8'h00;
		14'h2163:	ff_dbi <= 8'h00;
		14'h2164:	ff_dbi <= 8'h00;
		14'h2165:	ff_dbi <= 8'h00;
		14'h2166:	ff_dbi <= 8'h00;
		14'h2167:	ff_dbi <= 8'h00;
		14'h2168:	ff_dbi <= 8'h00;
		14'h2169:	ff_dbi <= 8'h00;
		14'h216a:	ff_dbi <= 8'h00;
		14'h216b:	ff_dbi <= 8'h00;
		14'h216c:	ff_dbi <= 8'h00;
		14'h216d:	ff_dbi <= 8'h00;
		14'h216e:	ff_dbi <= 8'h00;
		14'h216f:	ff_dbi <= 8'h00;
		14'h2170:	ff_dbi <= 8'h00;
		14'h2171:	ff_dbi <= 8'h00;
		14'h2172:	ff_dbi <= 8'h00;
		14'h2173:	ff_dbi <= 8'h00;
		14'h2174:	ff_dbi <= 8'h00;
		14'h2175:	ff_dbi <= 8'h00;
		14'h2176:	ff_dbi <= 8'h00;
		14'h2177:	ff_dbi <= 8'h00;
		14'h2178:	ff_dbi <= 8'h00;
		14'h2179:	ff_dbi <= 8'h00;
		14'h217a:	ff_dbi <= 8'h00;
		14'h217b:	ff_dbi <= 8'h00;
		14'h217c:	ff_dbi <= 8'h00;
		14'h217d:	ff_dbi <= 8'h00;
		14'h217e:	ff_dbi <= 8'h00;
		14'h217f:	ff_dbi <= 8'h00;
		14'h2180:	ff_dbi <= 8'h00;
		14'h2181:	ff_dbi <= 8'h00;
		14'h2182:	ff_dbi <= 8'h00;
		14'h2183:	ff_dbi <= 8'h00;
		14'h2184:	ff_dbi <= 8'h00;
		14'h2185:	ff_dbi <= 8'h00;
		14'h2186:	ff_dbi <= 8'h00;
		14'h2187:	ff_dbi <= 8'h00;
		14'h2188:	ff_dbi <= 8'h00;
		14'h2189:	ff_dbi <= 8'h00;
		14'h218a:	ff_dbi <= 8'h00;
		14'h218b:	ff_dbi <= 8'h00;
		14'h218c:	ff_dbi <= 8'h00;
		14'h218d:	ff_dbi <= 8'h00;
		14'h218e:	ff_dbi <= 8'h00;
		14'h218f:	ff_dbi <= 8'h00;
		14'h2190:	ff_dbi <= 8'h00;
		14'h2191:	ff_dbi <= 8'h00;
		14'h2192:	ff_dbi <= 8'h00;
		14'h2193:	ff_dbi <= 8'h00;
		14'h2194:	ff_dbi <= 8'h00;
		14'h2195:	ff_dbi <= 8'h00;
		14'h2196:	ff_dbi <= 8'h00;
		14'h2197:	ff_dbi <= 8'h00;
		14'h2198:	ff_dbi <= 8'h00;
		14'h2199:	ff_dbi <= 8'h00;
		14'h219a:	ff_dbi <= 8'h00;
		14'h219b:	ff_dbi <= 8'h00;
		14'h219c:	ff_dbi <= 8'h00;
		14'h219d:	ff_dbi <= 8'h00;
		14'h219e:	ff_dbi <= 8'h00;
		14'h219f:	ff_dbi <= 8'h00;
		14'h21a0:	ff_dbi <= 8'h00;
		14'h21a1:	ff_dbi <= 8'h00;
		14'h21a2:	ff_dbi <= 8'h00;
		14'h21a3:	ff_dbi <= 8'h00;
		14'h21a4:	ff_dbi <= 8'h00;
		14'h21a5:	ff_dbi <= 8'h00;
		14'h21a6:	ff_dbi <= 8'h00;
		14'h21a7:	ff_dbi <= 8'h00;
		14'h21a8:	ff_dbi <= 8'h00;
		14'h21a9:	ff_dbi <= 8'h00;
		14'h21aa:	ff_dbi <= 8'h00;
		14'h21ab:	ff_dbi <= 8'h00;
		14'h21ac:	ff_dbi <= 8'h00;
		14'h21ad:	ff_dbi <= 8'h00;
		14'h21ae:	ff_dbi <= 8'h00;
		14'h21af:	ff_dbi <= 8'h00;
		14'h21b0:	ff_dbi <= 8'h00;
		14'h21b1:	ff_dbi <= 8'h00;
		14'h21b2:	ff_dbi <= 8'h00;
		14'h21b3:	ff_dbi <= 8'h00;
		14'h21b4:	ff_dbi <= 8'h00;
		14'h21b5:	ff_dbi <= 8'h00;
		14'h21b6:	ff_dbi <= 8'h00;
		14'h21b7:	ff_dbi <= 8'h00;
		14'h21b8:	ff_dbi <= 8'h00;
		14'h21b9:	ff_dbi <= 8'h00;
		14'h21ba:	ff_dbi <= 8'h00;
		14'h21bb:	ff_dbi <= 8'h00;
		14'h21bc:	ff_dbi <= 8'h00;
		14'h21bd:	ff_dbi <= 8'h00;
		14'h21be:	ff_dbi <= 8'h00;
		14'h21bf:	ff_dbi <= 8'h00;
		14'h21c0:	ff_dbi <= 8'h00;
		14'h21c1:	ff_dbi <= 8'h00;
		14'h21c2:	ff_dbi <= 8'h00;
		14'h21c3:	ff_dbi <= 8'h00;
		14'h21c4:	ff_dbi <= 8'h00;
		14'h21c5:	ff_dbi <= 8'h00;
		14'h21c6:	ff_dbi <= 8'h00;
		14'h21c7:	ff_dbi <= 8'h00;
		14'h21c8:	ff_dbi <= 8'h00;
		14'h21c9:	ff_dbi <= 8'h00;
		14'h21ca:	ff_dbi <= 8'h00;
		14'h21cb:	ff_dbi <= 8'h00;
		14'h21cc:	ff_dbi <= 8'h00;
		14'h21cd:	ff_dbi <= 8'h00;
		14'h21ce:	ff_dbi <= 8'h00;
		14'h21cf:	ff_dbi <= 8'h00;
		14'h21d0:	ff_dbi <= 8'h00;
		14'h21d1:	ff_dbi <= 8'h00;
		14'h21d2:	ff_dbi <= 8'h00;
		14'h21d3:	ff_dbi <= 8'h00;
		14'h21d4:	ff_dbi <= 8'h00;
		14'h21d5:	ff_dbi <= 8'h00;
		14'h21d6:	ff_dbi <= 8'h00;
		14'h21d7:	ff_dbi <= 8'h00;
		14'h21d8:	ff_dbi <= 8'h00;
		14'h21d9:	ff_dbi <= 8'h00;
		14'h21da:	ff_dbi <= 8'h00;
		14'h21db:	ff_dbi <= 8'h00;
		14'h21dc:	ff_dbi <= 8'h00;
		14'h21dd:	ff_dbi <= 8'h00;
		14'h21de:	ff_dbi <= 8'h00;
		14'h21df:	ff_dbi <= 8'h00;
		14'h21e0:	ff_dbi <= 8'h00;
		14'h21e1:	ff_dbi <= 8'h00;
		14'h21e2:	ff_dbi <= 8'h00;
		14'h21e3:	ff_dbi <= 8'h00;
		14'h21e4:	ff_dbi <= 8'h00;
		14'h21e5:	ff_dbi <= 8'h00;
		14'h21e6:	ff_dbi <= 8'h00;
		14'h21e7:	ff_dbi <= 8'h00;
		14'h21e8:	ff_dbi <= 8'h00;
		14'h21e9:	ff_dbi <= 8'h00;
		14'h21ea:	ff_dbi <= 8'h00;
		14'h21eb:	ff_dbi <= 8'h00;
		14'h21ec:	ff_dbi <= 8'h00;
		14'h21ed:	ff_dbi <= 8'h00;
		14'h21ee:	ff_dbi <= 8'h00;
		14'h21ef:	ff_dbi <= 8'h00;
		14'h21f0:	ff_dbi <= 8'h00;
		14'h21f1:	ff_dbi <= 8'h00;
		14'h21f2:	ff_dbi <= 8'h00;
		14'h21f3:	ff_dbi <= 8'h00;
		14'h21f4:	ff_dbi <= 8'h00;
		14'h21f5:	ff_dbi <= 8'h00;
		14'h21f6:	ff_dbi <= 8'h00;
		14'h21f7:	ff_dbi <= 8'h00;
		14'h21f8:	ff_dbi <= 8'h00;
		14'h21f9:	ff_dbi <= 8'h00;
		14'h21fa:	ff_dbi <= 8'h00;
		14'h21fb:	ff_dbi <= 8'h00;
		14'h21fc:	ff_dbi <= 8'h00;
		14'h21fd:	ff_dbi <= 8'h00;
		14'h21fe:	ff_dbi <= 8'h00;
		14'h21ff:	ff_dbi <= 8'h00;
		14'h2200:	ff_dbi <= 8'h00;
		14'h2201:	ff_dbi <= 8'h00;
		14'h2202:	ff_dbi <= 8'h00;
		14'h2203:	ff_dbi <= 8'h00;
		14'h2204:	ff_dbi <= 8'h00;
		14'h2205:	ff_dbi <= 8'h00;
		14'h2206:	ff_dbi <= 8'h00;
		14'h2207:	ff_dbi <= 8'h00;
		14'h2208:	ff_dbi <= 8'h00;
		14'h2209:	ff_dbi <= 8'h00;
		14'h220a:	ff_dbi <= 8'h00;
		14'h220b:	ff_dbi <= 8'h00;
		14'h220c:	ff_dbi <= 8'h00;
		14'h220d:	ff_dbi <= 8'h00;
		14'h220e:	ff_dbi <= 8'h00;
		14'h220f:	ff_dbi <= 8'h00;
		14'h2210:	ff_dbi <= 8'h00;
		14'h2211:	ff_dbi <= 8'h00;
		14'h2212:	ff_dbi <= 8'h00;
		14'h2213:	ff_dbi <= 8'h00;
		14'h2214:	ff_dbi <= 8'h00;
		14'h2215:	ff_dbi <= 8'h00;
		14'h2216:	ff_dbi <= 8'h00;
		14'h2217:	ff_dbi <= 8'h00;
		14'h2218:	ff_dbi <= 8'h00;
		14'h2219:	ff_dbi <= 8'h00;
		14'h221a:	ff_dbi <= 8'h00;
		14'h221b:	ff_dbi <= 8'h00;
		14'h221c:	ff_dbi <= 8'h00;
		14'h221d:	ff_dbi <= 8'h00;
		14'h221e:	ff_dbi <= 8'h00;
		14'h221f:	ff_dbi <= 8'h00;
		14'h2220:	ff_dbi <= 8'h00;
		14'h2221:	ff_dbi <= 8'h00;
		14'h2222:	ff_dbi <= 8'h00;
		14'h2223:	ff_dbi <= 8'h00;
		14'h2224:	ff_dbi <= 8'h00;
		14'h2225:	ff_dbi <= 8'h00;
		14'h2226:	ff_dbi <= 8'h00;
		14'h2227:	ff_dbi <= 8'h00;
		14'h2228:	ff_dbi <= 8'h00;
		14'h2229:	ff_dbi <= 8'h00;
		14'h222a:	ff_dbi <= 8'h00;
		14'h222b:	ff_dbi <= 8'h00;
		14'h222c:	ff_dbi <= 8'h00;
		14'h222d:	ff_dbi <= 8'h00;
		14'h222e:	ff_dbi <= 8'h00;
		14'h222f:	ff_dbi <= 8'h00;
		14'h2230:	ff_dbi <= 8'h00;
		14'h2231:	ff_dbi <= 8'h00;
		14'h2232:	ff_dbi <= 8'h00;
		14'h2233:	ff_dbi <= 8'h00;
		14'h2234:	ff_dbi <= 8'h00;
		14'h2235:	ff_dbi <= 8'h00;
		14'h2236:	ff_dbi <= 8'h00;
		14'h2237:	ff_dbi <= 8'h00;
		14'h2238:	ff_dbi <= 8'h00;
		14'h2239:	ff_dbi <= 8'h00;
		14'h223a:	ff_dbi <= 8'h00;
		14'h223b:	ff_dbi <= 8'h00;
		14'h223c:	ff_dbi <= 8'h00;
		14'h223d:	ff_dbi <= 8'h00;
		14'h223e:	ff_dbi <= 8'h00;
		14'h223f:	ff_dbi <= 8'h00;
		14'h2240:	ff_dbi <= 8'h00;
		14'h2241:	ff_dbi <= 8'h00;
		14'h2242:	ff_dbi <= 8'h00;
		14'h2243:	ff_dbi <= 8'h00;
		14'h2244:	ff_dbi <= 8'h00;
		14'h2245:	ff_dbi <= 8'h00;
		14'h2246:	ff_dbi <= 8'h00;
		14'h2247:	ff_dbi <= 8'h00;
		14'h2248:	ff_dbi <= 8'h00;
		14'h2249:	ff_dbi <= 8'h00;
		14'h224a:	ff_dbi <= 8'h00;
		14'h224b:	ff_dbi <= 8'h00;
		14'h224c:	ff_dbi <= 8'h00;
		14'h224d:	ff_dbi <= 8'h00;
		14'h224e:	ff_dbi <= 8'h00;
		14'h224f:	ff_dbi <= 8'h00;
		14'h2250:	ff_dbi <= 8'h00;
		14'h2251:	ff_dbi <= 8'h00;
		14'h2252:	ff_dbi <= 8'h00;
		14'h2253:	ff_dbi <= 8'h00;
		14'h2254:	ff_dbi <= 8'h00;
		14'h2255:	ff_dbi <= 8'h00;
		14'h2256:	ff_dbi <= 8'h00;
		14'h2257:	ff_dbi <= 8'h00;
		14'h2258:	ff_dbi <= 8'h00;
		14'h2259:	ff_dbi <= 8'h00;
		14'h225a:	ff_dbi <= 8'h00;
		14'h225b:	ff_dbi <= 8'h00;
		14'h225c:	ff_dbi <= 8'h00;
		14'h225d:	ff_dbi <= 8'h00;
		14'h225e:	ff_dbi <= 8'h00;
		14'h225f:	ff_dbi <= 8'h00;
		14'h2260:	ff_dbi <= 8'h00;
		14'h2261:	ff_dbi <= 8'h00;
		14'h2262:	ff_dbi <= 8'h00;
		14'h2263:	ff_dbi <= 8'h00;
		14'h2264:	ff_dbi <= 8'h00;
		14'h2265:	ff_dbi <= 8'h00;
		14'h2266:	ff_dbi <= 8'h00;
		14'h2267:	ff_dbi <= 8'h00;
		14'h2268:	ff_dbi <= 8'h00;
		14'h2269:	ff_dbi <= 8'h00;
		14'h226a:	ff_dbi <= 8'h00;
		14'h226b:	ff_dbi <= 8'h00;
		14'h226c:	ff_dbi <= 8'h00;
		14'h226d:	ff_dbi <= 8'h00;
		14'h226e:	ff_dbi <= 8'h00;
		14'h226f:	ff_dbi <= 8'h00;
		14'h2270:	ff_dbi <= 8'h00;
		14'h2271:	ff_dbi <= 8'h00;
		14'h2272:	ff_dbi <= 8'h00;
		14'h2273:	ff_dbi <= 8'h00;
		14'h2274:	ff_dbi <= 8'h00;
		14'h2275:	ff_dbi <= 8'h00;
		14'h2276:	ff_dbi <= 8'h00;
		14'h2277:	ff_dbi <= 8'h00;
		14'h2278:	ff_dbi <= 8'h00;
		14'h2279:	ff_dbi <= 8'h00;
		14'h227a:	ff_dbi <= 8'h00;
		14'h227b:	ff_dbi <= 8'h00;
		14'h227c:	ff_dbi <= 8'h00;
		14'h227d:	ff_dbi <= 8'h00;
		14'h227e:	ff_dbi <= 8'h00;
		14'h227f:	ff_dbi <= 8'h00;
		14'h2280:	ff_dbi <= 8'h00;
		14'h2281:	ff_dbi <= 8'h00;
		14'h2282:	ff_dbi <= 8'h00;
		14'h2283:	ff_dbi <= 8'h00;
		14'h2284:	ff_dbi <= 8'h00;
		14'h2285:	ff_dbi <= 8'h00;
		14'h2286:	ff_dbi <= 8'h00;
		14'h2287:	ff_dbi <= 8'h00;
		14'h2288:	ff_dbi <= 8'h00;
		14'h2289:	ff_dbi <= 8'h00;
		14'h228a:	ff_dbi <= 8'h00;
		14'h228b:	ff_dbi <= 8'h00;
		14'h228c:	ff_dbi <= 8'h00;
		14'h228d:	ff_dbi <= 8'h00;
		14'h228e:	ff_dbi <= 8'h00;
		14'h228f:	ff_dbi <= 8'h00;
		14'h2290:	ff_dbi <= 8'h00;
		14'h2291:	ff_dbi <= 8'h00;
		14'h2292:	ff_dbi <= 8'h00;
		14'h2293:	ff_dbi <= 8'h00;
		14'h2294:	ff_dbi <= 8'h00;
		14'h2295:	ff_dbi <= 8'h00;
		14'h2296:	ff_dbi <= 8'h00;
		14'h2297:	ff_dbi <= 8'h00;
		14'h2298:	ff_dbi <= 8'h00;
		14'h2299:	ff_dbi <= 8'h00;
		14'h229a:	ff_dbi <= 8'h00;
		14'h229b:	ff_dbi <= 8'h00;
		14'h229c:	ff_dbi <= 8'h00;
		14'h229d:	ff_dbi <= 8'h00;
		14'h229e:	ff_dbi <= 8'h00;
		14'h229f:	ff_dbi <= 8'h00;
		14'h22a0:	ff_dbi <= 8'h00;
		14'h22a1:	ff_dbi <= 8'h00;
		14'h22a2:	ff_dbi <= 8'h00;
		14'h22a3:	ff_dbi <= 8'h00;
		14'h22a4:	ff_dbi <= 8'h00;
		14'h22a5:	ff_dbi <= 8'h00;
		14'h22a6:	ff_dbi <= 8'h00;
		14'h22a7:	ff_dbi <= 8'h00;
		14'h22a8:	ff_dbi <= 8'h00;
		14'h22a9:	ff_dbi <= 8'h00;
		14'h22aa:	ff_dbi <= 8'h00;
		14'h22ab:	ff_dbi <= 8'h00;
		14'h22ac:	ff_dbi <= 8'h00;
		14'h22ad:	ff_dbi <= 8'h00;
		14'h22ae:	ff_dbi <= 8'h00;
		14'h22af:	ff_dbi <= 8'h00;
		14'h22b0:	ff_dbi <= 8'h00;
		14'h22b1:	ff_dbi <= 8'h00;
		14'h22b2:	ff_dbi <= 8'h00;
		14'h22b3:	ff_dbi <= 8'h00;
		14'h22b4:	ff_dbi <= 8'h00;
		14'h22b5:	ff_dbi <= 8'h00;
		14'h22b6:	ff_dbi <= 8'h00;
		14'h22b7:	ff_dbi <= 8'h00;
		14'h22b8:	ff_dbi <= 8'h00;
		14'h22b9:	ff_dbi <= 8'h00;
		14'h22ba:	ff_dbi <= 8'h00;
		14'h22bb:	ff_dbi <= 8'h00;
		14'h22bc:	ff_dbi <= 8'h00;
		14'h22bd:	ff_dbi <= 8'h00;
		14'h22be:	ff_dbi <= 8'h00;
		14'h22bf:	ff_dbi <= 8'h00;
		14'h22c0:	ff_dbi <= 8'h00;
		14'h22c1:	ff_dbi <= 8'h00;
		14'h22c2:	ff_dbi <= 8'h00;
		14'h22c3:	ff_dbi <= 8'h00;
		14'h22c4:	ff_dbi <= 8'h00;
		14'h22c5:	ff_dbi <= 8'h00;
		14'h22c6:	ff_dbi <= 8'h00;
		14'h22c7:	ff_dbi <= 8'h00;
		14'h22c8:	ff_dbi <= 8'h00;
		14'h22c9:	ff_dbi <= 8'h00;
		14'h22ca:	ff_dbi <= 8'h00;
		14'h22cb:	ff_dbi <= 8'h00;
		14'h22cc:	ff_dbi <= 8'h00;
		14'h22cd:	ff_dbi <= 8'h00;
		14'h22ce:	ff_dbi <= 8'h00;
		14'h22cf:	ff_dbi <= 8'h00;
		14'h22d0:	ff_dbi <= 8'h00;
		14'h22d1:	ff_dbi <= 8'h00;
		14'h22d2:	ff_dbi <= 8'h00;
		14'h22d3:	ff_dbi <= 8'h00;
		14'h22d4:	ff_dbi <= 8'h00;
		14'h22d5:	ff_dbi <= 8'h00;
		14'h22d6:	ff_dbi <= 8'h00;
		14'h22d7:	ff_dbi <= 8'h00;
		14'h22d8:	ff_dbi <= 8'h00;
		14'h22d9:	ff_dbi <= 8'h00;
		14'h22da:	ff_dbi <= 8'h00;
		14'h22db:	ff_dbi <= 8'h00;
		14'h22dc:	ff_dbi <= 8'h00;
		14'h22dd:	ff_dbi <= 8'h00;
		14'h22de:	ff_dbi <= 8'h00;
		14'h22df:	ff_dbi <= 8'h00;
		14'h22e0:	ff_dbi <= 8'h00;
		14'h22e1:	ff_dbi <= 8'h00;
		14'h22e2:	ff_dbi <= 8'h00;
		14'h22e3:	ff_dbi <= 8'h00;
		14'h22e4:	ff_dbi <= 8'h00;
		14'h22e5:	ff_dbi <= 8'h00;
		14'h22e6:	ff_dbi <= 8'h00;
		14'h22e7:	ff_dbi <= 8'h00;
		14'h22e8:	ff_dbi <= 8'h00;
		14'h22e9:	ff_dbi <= 8'h00;
		14'h22ea:	ff_dbi <= 8'h00;
		14'h22eb:	ff_dbi <= 8'h00;
		14'h22ec:	ff_dbi <= 8'h00;
		14'h22ed:	ff_dbi <= 8'h00;
		14'h22ee:	ff_dbi <= 8'h00;
		14'h22ef:	ff_dbi <= 8'h00;
		14'h22f0:	ff_dbi <= 8'h00;
		14'h22f1:	ff_dbi <= 8'h00;
		14'h22f2:	ff_dbi <= 8'h00;
		14'h22f3:	ff_dbi <= 8'h00;
		14'h22f4:	ff_dbi <= 8'h00;
		14'h22f5:	ff_dbi <= 8'h00;
		14'h22f6:	ff_dbi <= 8'h00;
		14'h22f7:	ff_dbi <= 8'h00;
		14'h22f8:	ff_dbi <= 8'h00;
		14'h22f9:	ff_dbi <= 8'h00;
		14'h22fa:	ff_dbi <= 8'h00;
		14'h22fb:	ff_dbi <= 8'h00;
		14'h22fc:	ff_dbi <= 8'h00;
		14'h22fd:	ff_dbi <= 8'h00;
		14'h22fe:	ff_dbi <= 8'h00;
		14'h22ff:	ff_dbi <= 8'h00;
		14'h2300:	ff_dbi <= 8'h00;
		14'h2301:	ff_dbi <= 8'h00;
		14'h2302:	ff_dbi <= 8'h00;
		14'h2303:	ff_dbi <= 8'h00;
		14'h2304:	ff_dbi <= 8'h00;
		14'h2305:	ff_dbi <= 8'h00;
		14'h2306:	ff_dbi <= 8'h00;
		14'h2307:	ff_dbi <= 8'h00;
		14'h2308:	ff_dbi <= 8'h00;
		14'h2309:	ff_dbi <= 8'h00;
		14'h230a:	ff_dbi <= 8'h00;
		14'h230b:	ff_dbi <= 8'h00;
		14'h230c:	ff_dbi <= 8'h00;
		14'h230d:	ff_dbi <= 8'h00;
		14'h230e:	ff_dbi <= 8'h00;
		14'h230f:	ff_dbi <= 8'h00;
		14'h2310:	ff_dbi <= 8'h00;
		14'h2311:	ff_dbi <= 8'h00;
		14'h2312:	ff_dbi <= 8'h00;
		14'h2313:	ff_dbi <= 8'h00;
		14'h2314:	ff_dbi <= 8'h00;
		14'h2315:	ff_dbi <= 8'h00;
		14'h2316:	ff_dbi <= 8'h00;
		14'h2317:	ff_dbi <= 8'h00;
		14'h2318:	ff_dbi <= 8'h00;
		14'h2319:	ff_dbi <= 8'h00;
		14'h231a:	ff_dbi <= 8'h00;
		14'h231b:	ff_dbi <= 8'h00;
		14'h231c:	ff_dbi <= 8'h00;
		14'h231d:	ff_dbi <= 8'h00;
		14'h231e:	ff_dbi <= 8'h00;
		14'h231f:	ff_dbi <= 8'h00;
		14'h2320:	ff_dbi <= 8'h00;
		14'h2321:	ff_dbi <= 8'h00;
		14'h2322:	ff_dbi <= 8'h00;
		14'h2323:	ff_dbi <= 8'h00;
		14'h2324:	ff_dbi <= 8'h00;
		14'h2325:	ff_dbi <= 8'h00;
		14'h2326:	ff_dbi <= 8'h00;
		14'h2327:	ff_dbi <= 8'h00;
		14'h2328:	ff_dbi <= 8'h00;
		14'h2329:	ff_dbi <= 8'h00;
		14'h232a:	ff_dbi <= 8'h00;
		14'h232b:	ff_dbi <= 8'h00;
		14'h232c:	ff_dbi <= 8'h00;
		14'h232d:	ff_dbi <= 8'h00;
		14'h232e:	ff_dbi <= 8'h00;
		14'h232f:	ff_dbi <= 8'h00;
		14'h2330:	ff_dbi <= 8'h00;
		14'h2331:	ff_dbi <= 8'h00;
		14'h2332:	ff_dbi <= 8'h00;
		14'h2333:	ff_dbi <= 8'h00;
		14'h2334:	ff_dbi <= 8'h00;
		14'h2335:	ff_dbi <= 8'h00;
		14'h2336:	ff_dbi <= 8'h00;
		14'h2337:	ff_dbi <= 8'h00;
		14'h2338:	ff_dbi <= 8'h00;
		14'h2339:	ff_dbi <= 8'h00;
		14'h233a:	ff_dbi <= 8'h00;
		14'h233b:	ff_dbi <= 8'h00;
		14'h233c:	ff_dbi <= 8'h00;
		14'h233d:	ff_dbi <= 8'h00;
		14'h233e:	ff_dbi <= 8'h00;
		14'h233f:	ff_dbi <= 8'h00;
		14'h2340:	ff_dbi <= 8'h00;
		14'h2341:	ff_dbi <= 8'h00;
		14'h2342:	ff_dbi <= 8'h00;
		14'h2343:	ff_dbi <= 8'h00;
		14'h2344:	ff_dbi <= 8'h00;
		14'h2345:	ff_dbi <= 8'h00;
		14'h2346:	ff_dbi <= 8'h00;
		14'h2347:	ff_dbi <= 8'h00;
		14'h2348:	ff_dbi <= 8'h00;
		14'h2349:	ff_dbi <= 8'h00;
		14'h234a:	ff_dbi <= 8'h00;
		14'h234b:	ff_dbi <= 8'h00;
		14'h234c:	ff_dbi <= 8'h00;
		14'h234d:	ff_dbi <= 8'h00;
		14'h234e:	ff_dbi <= 8'h00;
		14'h234f:	ff_dbi <= 8'h00;
		14'h2350:	ff_dbi <= 8'h00;
		14'h2351:	ff_dbi <= 8'h00;
		14'h2352:	ff_dbi <= 8'h00;
		14'h2353:	ff_dbi <= 8'h00;
		14'h2354:	ff_dbi <= 8'h00;
		14'h2355:	ff_dbi <= 8'h00;
		14'h2356:	ff_dbi <= 8'h00;
		14'h2357:	ff_dbi <= 8'h00;
		14'h2358:	ff_dbi <= 8'h00;
		14'h2359:	ff_dbi <= 8'h00;
		14'h235a:	ff_dbi <= 8'h00;
		14'h235b:	ff_dbi <= 8'h00;
		14'h235c:	ff_dbi <= 8'h00;
		14'h235d:	ff_dbi <= 8'h00;
		14'h235e:	ff_dbi <= 8'h00;
		14'h235f:	ff_dbi <= 8'h00;
		14'h2360:	ff_dbi <= 8'h00;
		14'h2361:	ff_dbi <= 8'h00;
		14'h2362:	ff_dbi <= 8'h00;
		14'h2363:	ff_dbi <= 8'h00;
		14'h2364:	ff_dbi <= 8'h00;
		14'h2365:	ff_dbi <= 8'h00;
		14'h2366:	ff_dbi <= 8'h00;
		14'h2367:	ff_dbi <= 8'h00;
		14'h2368:	ff_dbi <= 8'h00;
		14'h2369:	ff_dbi <= 8'h00;
		14'h236a:	ff_dbi <= 8'h00;
		14'h236b:	ff_dbi <= 8'h00;
		14'h236c:	ff_dbi <= 8'h00;
		14'h236d:	ff_dbi <= 8'h00;
		14'h236e:	ff_dbi <= 8'h00;
		14'h236f:	ff_dbi <= 8'h00;
		14'h2370:	ff_dbi <= 8'h00;
		14'h2371:	ff_dbi <= 8'h00;
		14'h2372:	ff_dbi <= 8'h00;
		14'h2373:	ff_dbi <= 8'h00;
		14'h2374:	ff_dbi <= 8'h00;
		14'h2375:	ff_dbi <= 8'h00;
		14'h2376:	ff_dbi <= 8'h00;
		14'h2377:	ff_dbi <= 8'h00;
		14'h2378:	ff_dbi <= 8'h00;
		14'h2379:	ff_dbi <= 8'h00;
		14'h237a:	ff_dbi <= 8'h00;
		14'h237b:	ff_dbi <= 8'h00;
		14'h237c:	ff_dbi <= 8'h00;
		14'h237d:	ff_dbi <= 8'h00;
		14'h237e:	ff_dbi <= 8'h00;
		14'h237f:	ff_dbi <= 8'h00;
		14'h2380:	ff_dbi <= 8'h00;
		14'h2381:	ff_dbi <= 8'h00;
		14'h2382:	ff_dbi <= 8'h00;
		14'h2383:	ff_dbi <= 8'h00;
		14'h2384:	ff_dbi <= 8'h00;
		14'h2385:	ff_dbi <= 8'h00;
		14'h2386:	ff_dbi <= 8'h00;
		14'h2387:	ff_dbi <= 8'h00;
		14'h2388:	ff_dbi <= 8'h00;
		14'h2389:	ff_dbi <= 8'h00;
		14'h238a:	ff_dbi <= 8'h00;
		14'h238b:	ff_dbi <= 8'h00;
		14'h238c:	ff_dbi <= 8'h00;
		14'h238d:	ff_dbi <= 8'h00;
		14'h238e:	ff_dbi <= 8'h00;
		14'h238f:	ff_dbi <= 8'h00;
		14'h2390:	ff_dbi <= 8'h00;
		14'h2391:	ff_dbi <= 8'h00;
		14'h2392:	ff_dbi <= 8'h00;
		14'h2393:	ff_dbi <= 8'h00;
		14'h2394:	ff_dbi <= 8'h00;
		14'h2395:	ff_dbi <= 8'h00;
		14'h2396:	ff_dbi <= 8'h00;
		14'h2397:	ff_dbi <= 8'h00;
		14'h2398:	ff_dbi <= 8'h00;
		14'h2399:	ff_dbi <= 8'h00;
		14'h239a:	ff_dbi <= 8'h00;
		14'h239b:	ff_dbi <= 8'h00;
		14'h239c:	ff_dbi <= 8'h00;
		14'h239d:	ff_dbi <= 8'h00;
		14'h239e:	ff_dbi <= 8'h00;
		14'h239f:	ff_dbi <= 8'h00;
		14'h23a0:	ff_dbi <= 8'h00;
		14'h23a1:	ff_dbi <= 8'h00;
		14'h23a2:	ff_dbi <= 8'h00;
		14'h23a3:	ff_dbi <= 8'h00;
		14'h23a4:	ff_dbi <= 8'h00;
		14'h23a5:	ff_dbi <= 8'h00;
		14'h23a6:	ff_dbi <= 8'h00;
		14'h23a7:	ff_dbi <= 8'h00;
		14'h23a8:	ff_dbi <= 8'h00;
		14'h23a9:	ff_dbi <= 8'h00;
		14'h23aa:	ff_dbi <= 8'h00;
		14'h23ab:	ff_dbi <= 8'h00;
		14'h23ac:	ff_dbi <= 8'h00;
		14'h23ad:	ff_dbi <= 8'h00;
		14'h23ae:	ff_dbi <= 8'h00;
		14'h23af:	ff_dbi <= 8'h00;
		14'h23b0:	ff_dbi <= 8'h00;
		14'h23b1:	ff_dbi <= 8'h00;
		14'h23b2:	ff_dbi <= 8'h00;
		14'h23b3:	ff_dbi <= 8'h00;
		14'h23b4:	ff_dbi <= 8'h00;
		14'h23b5:	ff_dbi <= 8'h00;
		14'h23b6:	ff_dbi <= 8'h00;
		14'h23b7:	ff_dbi <= 8'h00;
		14'h23b8:	ff_dbi <= 8'h00;
		14'h23b9:	ff_dbi <= 8'h00;
		14'h23ba:	ff_dbi <= 8'h00;
		14'h23bb:	ff_dbi <= 8'h00;
		14'h23bc:	ff_dbi <= 8'h00;
		14'h23bd:	ff_dbi <= 8'h00;
		14'h23be:	ff_dbi <= 8'h00;
		14'h23bf:	ff_dbi <= 8'h00;
		14'h23c0:	ff_dbi <= 8'h00;
		14'h23c1:	ff_dbi <= 8'h00;
		14'h23c2:	ff_dbi <= 8'h00;
		14'h23c3:	ff_dbi <= 8'h00;
		14'h23c4:	ff_dbi <= 8'h00;
		14'h23c5:	ff_dbi <= 8'h00;
		14'h23c6:	ff_dbi <= 8'h00;
		14'h23c7:	ff_dbi <= 8'h00;
		14'h23c8:	ff_dbi <= 8'h00;
		14'h23c9:	ff_dbi <= 8'h00;
		14'h23ca:	ff_dbi <= 8'h00;
		14'h23cb:	ff_dbi <= 8'h00;
		14'h23cc:	ff_dbi <= 8'h00;
		14'h23cd:	ff_dbi <= 8'h00;
		14'h23ce:	ff_dbi <= 8'h00;
		14'h23cf:	ff_dbi <= 8'h00;
		14'h23d0:	ff_dbi <= 8'h00;
		14'h23d1:	ff_dbi <= 8'h00;
		14'h23d2:	ff_dbi <= 8'h00;
		14'h23d3:	ff_dbi <= 8'h00;
		14'h23d4:	ff_dbi <= 8'h00;
		14'h23d5:	ff_dbi <= 8'h00;
		14'h23d6:	ff_dbi <= 8'h00;
		14'h23d7:	ff_dbi <= 8'h00;
		14'h23d8:	ff_dbi <= 8'h00;
		14'h23d9:	ff_dbi <= 8'h00;
		14'h23da:	ff_dbi <= 8'h00;
		14'h23db:	ff_dbi <= 8'h00;
		14'h23dc:	ff_dbi <= 8'h00;
		14'h23dd:	ff_dbi <= 8'h00;
		14'h23de:	ff_dbi <= 8'h00;
		14'h23df:	ff_dbi <= 8'h00;
		14'h23e0:	ff_dbi <= 8'h00;
		14'h23e1:	ff_dbi <= 8'h00;
		14'h23e2:	ff_dbi <= 8'h00;
		14'h23e3:	ff_dbi <= 8'h00;
		14'h23e4:	ff_dbi <= 8'h00;
		14'h23e5:	ff_dbi <= 8'h00;
		14'h23e6:	ff_dbi <= 8'h00;
		14'h23e7:	ff_dbi <= 8'h00;
		14'h23e8:	ff_dbi <= 8'h00;
		14'h23e9:	ff_dbi <= 8'h00;
		14'h23ea:	ff_dbi <= 8'h00;
		14'h23eb:	ff_dbi <= 8'h00;
		14'h23ec:	ff_dbi <= 8'h00;
		14'h23ed:	ff_dbi <= 8'h00;
		14'h23ee:	ff_dbi <= 8'h00;
		14'h23ef:	ff_dbi <= 8'h00;
		14'h23f0:	ff_dbi <= 8'h00;
		14'h23f1:	ff_dbi <= 8'h00;
		14'h23f2:	ff_dbi <= 8'h00;
		14'h23f3:	ff_dbi <= 8'h00;
		14'h23f4:	ff_dbi <= 8'h00;
		14'h23f5:	ff_dbi <= 8'h00;
		14'h23f6:	ff_dbi <= 8'h00;
		14'h23f7:	ff_dbi <= 8'h00;
		14'h23f8:	ff_dbi <= 8'h00;
		14'h23f9:	ff_dbi <= 8'h00;
		14'h23fa:	ff_dbi <= 8'h00;
		14'h23fb:	ff_dbi <= 8'h00;
		14'h23fc:	ff_dbi <= 8'h00;
		14'h23fd:	ff_dbi <= 8'h00;
		14'h23fe:	ff_dbi <= 8'h00;
		14'h23ff:	ff_dbi <= 8'h00;
		14'h2400:	ff_dbi <= 8'h00;
		14'h2401:	ff_dbi <= 8'h00;
		14'h2402:	ff_dbi <= 8'h00;
		14'h2403:	ff_dbi <= 8'h00;
		14'h2404:	ff_dbi <= 8'h00;
		14'h2405:	ff_dbi <= 8'h00;
		14'h2406:	ff_dbi <= 8'h00;
		14'h2407:	ff_dbi <= 8'h00;
		14'h2408:	ff_dbi <= 8'h00;
		14'h2409:	ff_dbi <= 8'h00;
		14'h240a:	ff_dbi <= 8'h00;
		14'h240b:	ff_dbi <= 8'h00;
		14'h240c:	ff_dbi <= 8'h00;
		14'h240d:	ff_dbi <= 8'h00;
		14'h240e:	ff_dbi <= 8'h00;
		14'h240f:	ff_dbi <= 8'h00;
		14'h2410:	ff_dbi <= 8'h00;
		14'h2411:	ff_dbi <= 8'h00;
		14'h2412:	ff_dbi <= 8'h00;
		14'h2413:	ff_dbi <= 8'h00;
		14'h2414:	ff_dbi <= 8'h00;
		14'h2415:	ff_dbi <= 8'h00;
		14'h2416:	ff_dbi <= 8'h00;
		14'h2417:	ff_dbi <= 8'h00;
		14'h2418:	ff_dbi <= 8'h00;
		14'h2419:	ff_dbi <= 8'h00;
		14'h241a:	ff_dbi <= 8'h00;
		14'h241b:	ff_dbi <= 8'h00;
		14'h241c:	ff_dbi <= 8'h00;
		14'h241d:	ff_dbi <= 8'h00;
		14'h241e:	ff_dbi <= 8'h00;
		14'h241f:	ff_dbi <= 8'h00;
		14'h2420:	ff_dbi <= 8'h00;
		14'h2421:	ff_dbi <= 8'h00;
		14'h2422:	ff_dbi <= 8'h00;
		14'h2423:	ff_dbi <= 8'h00;
		14'h2424:	ff_dbi <= 8'h00;
		14'h2425:	ff_dbi <= 8'h00;
		14'h2426:	ff_dbi <= 8'h00;
		14'h2427:	ff_dbi <= 8'h00;
		14'h2428:	ff_dbi <= 8'h00;
		14'h2429:	ff_dbi <= 8'h00;
		14'h242a:	ff_dbi <= 8'h00;
		14'h242b:	ff_dbi <= 8'h00;
		14'h242c:	ff_dbi <= 8'h00;
		14'h242d:	ff_dbi <= 8'h00;
		14'h242e:	ff_dbi <= 8'h00;
		14'h242f:	ff_dbi <= 8'h00;
		14'h2430:	ff_dbi <= 8'h00;
		14'h2431:	ff_dbi <= 8'h00;
		14'h2432:	ff_dbi <= 8'h00;
		14'h2433:	ff_dbi <= 8'h00;
		14'h2434:	ff_dbi <= 8'h00;
		14'h2435:	ff_dbi <= 8'h00;
		14'h2436:	ff_dbi <= 8'h00;
		14'h2437:	ff_dbi <= 8'h00;
		14'h2438:	ff_dbi <= 8'h00;
		14'h2439:	ff_dbi <= 8'h00;
		14'h243a:	ff_dbi <= 8'h00;
		14'h243b:	ff_dbi <= 8'h00;
		14'h243c:	ff_dbi <= 8'h00;
		14'h243d:	ff_dbi <= 8'h00;
		14'h243e:	ff_dbi <= 8'h00;
		14'h243f:	ff_dbi <= 8'h00;
		14'h2440:	ff_dbi <= 8'h00;
		14'h2441:	ff_dbi <= 8'h00;
		14'h2442:	ff_dbi <= 8'h00;
		14'h2443:	ff_dbi <= 8'h00;
		14'h2444:	ff_dbi <= 8'h00;
		14'h2445:	ff_dbi <= 8'h00;
		14'h2446:	ff_dbi <= 8'h00;
		14'h2447:	ff_dbi <= 8'h00;
		14'h2448:	ff_dbi <= 8'h00;
		14'h2449:	ff_dbi <= 8'h00;
		14'h244a:	ff_dbi <= 8'h00;
		14'h244b:	ff_dbi <= 8'h00;
		14'h244c:	ff_dbi <= 8'h00;
		14'h244d:	ff_dbi <= 8'h00;
		14'h244e:	ff_dbi <= 8'h00;
		14'h244f:	ff_dbi <= 8'h00;
		14'h2450:	ff_dbi <= 8'h00;
		14'h2451:	ff_dbi <= 8'h00;
		14'h2452:	ff_dbi <= 8'h00;
		14'h2453:	ff_dbi <= 8'h00;
		14'h2454:	ff_dbi <= 8'h00;
		14'h2455:	ff_dbi <= 8'h00;
		14'h2456:	ff_dbi <= 8'h00;
		14'h2457:	ff_dbi <= 8'h00;
		14'h2458:	ff_dbi <= 8'h00;
		14'h2459:	ff_dbi <= 8'h00;
		14'h245a:	ff_dbi <= 8'h00;
		14'h245b:	ff_dbi <= 8'h00;
		14'h245c:	ff_dbi <= 8'h00;
		14'h245d:	ff_dbi <= 8'h00;
		14'h245e:	ff_dbi <= 8'h00;
		14'h245f:	ff_dbi <= 8'h00;
		14'h2460:	ff_dbi <= 8'h00;
		14'h2461:	ff_dbi <= 8'h00;
		14'h2462:	ff_dbi <= 8'h00;
		14'h2463:	ff_dbi <= 8'h00;
		14'h2464:	ff_dbi <= 8'h00;
		14'h2465:	ff_dbi <= 8'h00;
		14'h2466:	ff_dbi <= 8'h00;
		14'h2467:	ff_dbi <= 8'h00;
		14'h2468:	ff_dbi <= 8'h00;
		14'h2469:	ff_dbi <= 8'h00;
		14'h246a:	ff_dbi <= 8'h00;
		14'h246b:	ff_dbi <= 8'h00;
		14'h246c:	ff_dbi <= 8'h00;
		14'h246d:	ff_dbi <= 8'h00;
		14'h246e:	ff_dbi <= 8'h00;
		14'h246f:	ff_dbi <= 8'h00;
		14'h2470:	ff_dbi <= 8'h00;
		14'h2471:	ff_dbi <= 8'h00;
		14'h2472:	ff_dbi <= 8'h00;
		14'h2473:	ff_dbi <= 8'h00;
		14'h2474:	ff_dbi <= 8'h00;
		14'h2475:	ff_dbi <= 8'h00;
		14'h2476:	ff_dbi <= 8'h00;
		14'h2477:	ff_dbi <= 8'h00;
		14'h2478:	ff_dbi <= 8'h00;
		14'h2479:	ff_dbi <= 8'h00;
		14'h247a:	ff_dbi <= 8'h00;
		14'h247b:	ff_dbi <= 8'h00;
		14'h247c:	ff_dbi <= 8'h00;
		14'h247d:	ff_dbi <= 8'h00;
		14'h247e:	ff_dbi <= 8'h00;
		14'h247f:	ff_dbi <= 8'h00;
		14'h2480:	ff_dbi <= 8'h00;
		14'h2481:	ff_dbi <= 8'h00;
		14'h2482:	ff_dbi <= 8'h00;
		14'h2483:	ff_dbi <= 8'h00;
		14'h2484:	ff_dbi <= 8'h00;
		14'h2485:	ff_dbi <= 8'h00;
		14'h2486:	ff_dbi <= 8'h00;
		14'h2487:	ff_dbi <= 8'h00;
		14'h2488:	ff_dbi <= 8'h00;
		14'h2489:	ff_dbi <= 8'h00;
		14'h248a:	ff_dbi <= 8'h00;
		14'h248b:	ff_dbi <= 8'h00;
		14'h248c:	ff_dbi <= 8'h00;
		14'h248d:	ff_dbi <= 8'h00;
		14'h248e:	ff_dbi <= 8'h00;
		14'h248f:	ff_dbi <= 8'h00;
		14'h2490:	ff_dbi <= 8'h00;
		14'h2491:	ff_dbi <= 8'h00;
		14'h2492:	ff_dbi <= 8'h00;
		14'h2493:	ff_dbi <= 8'h00;
		14'h2494:	ff_dbi <= 8'h00;
		14'h2495:	ff_dbi <= 8'h00;
		14'h2496:	ff_dbi <= 8'h00;
		14'h2497:	ff_dbi <= 8'h00;
		14'h2498:	ff_dbi <= 8'h00;
		14'h2499:	ff_dbi <= 8'h00;
		14'h249a:	ff_dbi <= 8'h00;
		14'h249b:	ff_dbi <= 8'h00;
		14'h249c:	ff_dbi <= 8'h00;
		14'h249d:	ff_dbi <= 8'h00;
		14'h249e:	ff_dbi <= 8'h00;
		14'h249f:	ff_dbi <= 8'h00;
		14'h24a0:	ff_dbi <= 8'h00;
		14'h24a1:	ff_dbi <= 8'h00;
		14'h24a2:	ff_dbi <= 8'h00;
		14'h24a3:	ff_dbi <= 8'h00;
		14'h24a4:	ff_dbi <= 8'h00;
		14'h24a5:	ff_dbi <= 8'h00;
		14'h24a6:	ff_dbi <= 8'h00;
		14'h24a7:	ff_dbi <= 8'h00;
		14'h24a8:	ff_dbi <= 8'h00;
		14'h24a9:	ff_dbi <= 8'h00;
		14'h24aa:	ff_dbi <= 8'h00;
		14'h24ab:	ff_dbi <= 8'h00;
		14'h24ac:	ff_dbi <= 8'h00;
		14'h24ad:	ff_dbi <= 8'h00;
		14'h24ae:	ff_dbi <= 8'h00;
		14'h24af:	ff_dbi <= 8'h00;
		14'h24b0:	ff_dbi <= 8'h00;
		14'h24b1:	ff_dbi <= 8'h00;
		14'h24b2:	ff_dbi <= 8'h00;
		14'h24b3:	ff_dbi <= 8'h00;
		14'h24b4:	ff_dbi <= 8'h00;
		14'h24b5:	ff_dbi <= 8'h00;
		14'h24b6:	ff_dbi <= 8'h00;
		14'h24b7:	ff_dbi <= 8'h00;
		14'h24b8:	ff_dbi <= 8'h00;
		14'h24b9:	ff_dbi <= 8'h00;
		14'h24ba:	ff_dbi <= 8'h00;
		14'h24bb:	ff_dbi <= 8'h00;
		14'h24bc:	ff_dbi <= 8'h00;
		14'h24bd:	ff_dbi <= 8'h00;
		14'h24be:	ff_dbi <= 8'h00;
		14'h24bf:	ff_dbi <= 8'h00;
		14'h24c0:	ff_dbi <= 8'h00;
		14'h24c1:	ff_dbi <= 8'h00;
		14'h24c2:	ff_dbi <= 8'h00;
		14'h24c3:	ff_dbi <= 8'h00;
		14'h24c4:	ff_dbi <= 8'h00;
		14'h24c5:	ff_dbi <= 8'h00;
		14'h24c6:	ff_dbi <= 8'h00;
		14'h24c7:	ff_dbi <= 8'h00;
		14'h24c8:	ff_dbi <= 8'h00;
		14'h24c9:	ff_dbi <= 8'h00;
		14'h24ca:	ff_dbi <= 8'h00;
		14'h24cb:	ff_dbi <= 8'h00;
		14'h24cc:	ff_dbi <= 8'h00;
		14'h24cd:	ff_dbi <= 8'h00;
		14'h24ce:	ff_dbi <= 8'h00;
		14'h24cf:	ff_dbi <= 8'h00;
		14'h24d0:	ff_dbi <= 8'h00;
		14'h24d1:	ff_dbi <= 8'h00;
		14'h24d2:	ff_dbi <= 8'h00;
		14'h24d3:	ff_dbi <= 8'h00;
		14'h24d4:	ff_dbi <= 8'h00;
		14'h24d5:	ff_dbi <= 8'h00;
		14'h24d6:	ff_dbi <= 8'h00;
		14'h24d7:	ff_dbi <= 8'h00;
		14'h24d8:	ff_dbi <= 8'h00;
		14'h24d9:	ff_dbi <= 8'h00;
		14'h24da:	ff_dbi <= 8'h00;
		14'h24db:	ff_dbi <= 8'h00;
		14'h24dc:	ff_dbi <= 8'h00;
		14'h24dd:	ff_dbi <= 8'h00;
		14'h24de:	ff_dbi <= 8'h00;
		14'h24df:	ff_dbi <= 8'h00;
		14'h24e0:	ff_dbi <= 8'h00;
		14'h24e1:	ff_dbi <= 8'h00;
		14'h24e2:	ff_dbi <= 8'h00;
		14'h24e3:	ff_dbi <= 8'h00;
		14'h24e4:	ff_dbi <= 8'h00;
		14'h24e5:	ff_dbi <= 8'h00;
		14'h24e6:	ff_dbi <= 8'h00;
		14'h24e7:	ff_dbi <= 8'h00;
		14'h24e8:	ff_dbi <= 8'h00;
		14'h24e9:	ff_dbi <= 8'h00;
		14'h24ea:	ff_dbi <= 8'h00;
		14'h24eb:	ff_dbi <= 8'h00;
		14'h24ec:	ff_dbi <= 8'h00;
		14'h24ed:	ff_dbi <= 8'h00;
		14'h24ee:	ff_dbi <= 8'h00;
		14'h24ef:	ff_dbi <= 8'h00;
		14'h24f0:	ff_dbi <= 8'h00;
		14'h24f1:	ff_dbi <= 8'h00;
		14'h24f2:	ff_dbi <= 8'h00;
		14'h24f3:	ff_dbi <= 8'h00;
		14'h24f4:	ff_dbi <= 8'h00;
		14'h24f5:	ff_dbi <= 8'h00;
		14'h24f6:	ff_dbi <= 8'h00;
		14'h24f7:	ff_dbi <= 8'h00;
		14'h24f8:	ff_dbi <= 8'h00;
		14'h24f9:	ff_dbi <= 8'h00;
		14'h24fa:	ff_dbi <= 8'h00;
		14'h24fb:	ff_dbi <= 8'h00;
		14'h24fc:	ff_dbi <= 8'h00;
		14'h24fd:	ff_dbi <= 8'h00;
		14'h24fe:	ff_dbi <= 8'h00;
		14'h24ff:	ff_dbi <= 8'h00;
		14'h2500:	ff_dbi <= 8'h00;
		14'h2501:	ff_dbi <= 8'h00;
		14'h2502:	ff_dbi <= 8'h00;
		14'h2503:	ff_dbi <= 8'h00;
		14'h2504:	ff_dbi <= 8'h00;
		14'h2505:	ff_dbi <= 8'h00;
		14'h2506:	ff_dbi <= 8'h00;
		14'h2507:	ff_dbi <= 8'h00;
		14'h2508:	ff_dbi <= 8'h00;
		14'h2509:	ff_dbi <= 8'h00;
		14'h250a:	ff_dbi <= 8'h00;
		14'h250b:	ff_dbi <= 8'h00;
		14'h250c:	ff_dbi <= 8'h00;
		14'h250d:	ff_dbi <= 8'h00;
		14'h250e:	ff_dbi <= 8'h00;
		14'h250f:	ff_dbi <= 8'h00;
		14'h2510:	ff_dbi <= 8'h00;
		14'h2511:	ff_dbi <= 8'h00;
		14'h2512:	ff_dbi <= 8'h00;
		14'h2513:	ff_dbi <= 8'h00;
		14'h2514:	ff_dbi <= 8'h00;
		14'h2515:	ff_dbi <= 8'h00;
		14'h2516:	ff_dbi <= 8'h00;
		14'h2517:	ff_dbi <= 8'h00;
		14'h2518:	ff_dbi <= 8'h00;
		14'h2519:	ff_dbi <= 8'h00;
		14'h251a:	ff_dbi <= 8'h00;
		14'h251b:	ff_dbi <= 8'h00;
		14'h251c:	ff_dbi <= 8'h00;
		14'h251d:	ff_dbi <= 8'h00;
		14'h251e:	ff_dbi <= 8'h00;
		14'h251f:	ff_dbi <= 8'h00;
		14'h2520:	ff_dbi <= 8'h00;
		14'h2521:	ff_dbi <= 8'h00;
		14'h2522:	ff_dbi <= 8'h00;
		14'h2523:	ff_dbi <= 8'h00;
		14'h2524:	ff_dbi <= 8'h00;
		14'h2525:	ff_dbi <= 8'h00;
		14'h2526:	ff_dbi <= 8'h00;
		14'h2527:	ff_dbi <= 8'h00;
		14'h2528:	ff_dbi <= 8'h00;
		14'h2529:	ff_dbi <= 8'h00;
		14'h252a:	ff_dbi <= 8'h00;
		14'h252b:	ff_dbi <= 8'h00;
		14'h252c:	ff_dbi <= 8'h00;
		14'h252d:	ff_dbi <= 8'h00;
		14'h252e:	ff_dbi <= 8'h00;
		14'h252f:	ff_dbi <= 8'h00;
		14'h2530:	ff_dbi <= 8'h00;
		14'h2531:	ff_dbi <= 8'h00;
		14'h2532:	ff_dbi <= 8'h00;
		14'h2533:	ff_dbi <= 8'h00;
		14'h2534:	ff_dbi <= 8'h00;
		14'h2535:	ff_dbi <= 8'h00;
		14'h2536:	ff_dbi <= 8'h00;
		14'h2537:	ff_dbi <= 8'h00;
		14'h2538:	ff_dbi <= 8'h00;
		14'h2539:	ff_dbi <= 8'h00;
		14'h253a:	ff_dbi <= 8'h00;
		14'h253b:	ff_dbi <= 8'h00;
		14'h253c:	ff_dbi <= 8'h00;
		14'h253d:	ff_dbi <= 8'h00;
		14'h253e:	ff_dbi <= 8'h00;
		14'h253f:	ff_dbi <= 8'h00;
		14'h2540:	ff_dbi <= 8'h00;
		14'h2541:	ff_dbi <= 8'h00;
		14'h2542:	ff_dbi <= 8'h00;
		14'h2543:	ff_dbi <= 8'h00;
		14'h2544:	ff_dbi <= 8'h00;
		14'h2545:	ff_dbi <= 8'h00;
		14'h2546:	ff_dbi <= 8'h00;
		14'h2547:	ff_dbi <= 8'h00;
		14'h2548:	ff_dbi <= 8'h00;
		14'h2549:	ff_dbi <= 8'h00;
		14'h254a:	ff_dbi <= 8'h00;
		14'h254b:	ff_dbi <= 8'h00;
		14'h254c:	ff_dbi <= 8'h00;
		14'h254d:	ff_dbi <= 8'h00;
		14'h254e:	ff_dbi <= 8'h00;
		14'h254f:	ff_dbi <= 8'h00;
		14'h2550:	ff_dbi <= 8'h00;
		14'h2551:	ff_dbi <= 8'h00;
		14'h2552:	ff_dbi <= 8'h00;
		14'h2553:	ff_dbi <= 8'h00;
		14'h2554:	ff_dbi <= 8'h00;
		14'h2555:	ff_dbi <= 8'h00;
		14'h2556:	ff_dbi <= 8'h00;
		14'h2557:	ff_dbi <= 8'h00;
		14'h2558:	ff_dbi <= 8'h00;
		14'h2559:	ff_dbi <= 8'h00;
		14'h255a:	ff_dbi <= 8'h00;
		14'h255b:	ff_dbi <= 8'h00;
		14'h255c:	ff_dbi <= 8'h00;
		14'h255d:	ff_dbi <= 8'h00;
		14'h255e:	ff_dbi <= 8'h00;
		14'h255f:	ff_dbi <= 8'h00;
		14'h2560:	ff_dbi <= 8'h00;
		14'h2561:	ff_dbi <= 8'h00;
		14'h2562:	ff_dbi <= 8'h00;
		14'h2563:	ff_dbi <= 8'h00;
		14'h2564:	ff_dbi <= 8'h00;
		14'h2565:	ff_dbi <= 8'h00;
		14'h2566:	ff_dbi <= 8'h00;
		14'h2567:	ff_dbi <= 8'h00;
		14'h2568:	ff_dbi <= 8'h00;
		14'h2569:	ff_dbi <= 8'h00;
		14'h256a:	ff_dbi <= 8'h00;
		14'h256b:	ff_dbi <= 8'h00;
		14'h256c:	ff_dbi <= 8'h00;
		14'h256d:	ff_dbi <= 8'h00;
		14'h256e:	ff_dbi <= 8'h00;
		14'h256f:	ff_dbi <= 8'h00;
		14'h2570:	ff_dbi <= 8'h00;
		14'h2571:	ff_dbi <= 8'h00;
		14'h2572:	ff_dbi <= 8'h00;
		14'h2573:	ff_dbi <= 8'h00;
		14'h2574:	ff_dbi <= 8'h00;
		14'h2575:	ff_dbi <= 8'h00;
		14'h2576:	ff_dbi <= 8'h00;
		14'h2577:	ff_dbi <= 8'h00;
		14'h2578:	ff_dbi <= 8'h00;
		14'h2579:	ff_dbi <= 8'h00;
		14'h257a:	ff_dbi <= 8'h00;
		14'h257b:	ff_dbi <= 8'h00;
		14'h257c:	ff_dbi <= 8'h00;
		14'h257d:	ff_dbi <= 8'h00;
		14'h257e:	ff_dbi <= 8'h00;
		14'h257f:	ff_dbi <= 8'h00;
		14'h2580:	ff_dbi <= 8'h00;
		14'h2581:	ff_dbi <= 8'h00;
		14'h2582:	ff_dbi <= 8'h00;
		14'h2583:	ff_dbi <= 8'h00;
		14'h2584:	ff_dbi <= 8'h00;
		14'h2585:	ff_dbi <= 8'h00;
		14'h2586:	ff_dbi <= 8'h00;
		14'h2587:	ff_dbi <= 8'h00;
		14'h2588:	ff_dbi <= 8'h00;
		14'h2589:	ff_dbi <= 8'h00;
		14'h258a:	ff_dbi <= 8'h00;
		14'h258b:	ff_dbi <= 8'h00;
		14'h258c:	ff_dbi <= 8'h00;
		14'h258d:	ff_dbi <= 8'h00;
		14'h258e:	ff_dbi <= 8'h00;
		14'h258f:	ff_dbi <= 8'h00;
		14'h2590:	ff_dbi <= 8'h00;
		14'h2591:	ff_dbi <= 8'h00;
		14'h2592:	ff_dbi <= 8'h00;
		14'h2593:	ff_dbi <= 8'h00;
		14'h2594:	ff_dbi <= 8'h00;
		14'h2595:	ff_dbi <= 8'h00;
		14'h2596:	ff_dbi <= 8'h00;
		14'h2597:	ff_dbi <= 8'h00;
		14'h2598:	ff_dbi <= 8'h00;
		14'h2599:	ff_dbi <= 8'h00;
		14'h259a:	ff_dbi <= 8'h00;
		14'h259b:	ff_dbi <= 8'h00;
		14'h259c:	ff_dbi <= 8'h00;
		14'h259d:	ff_dbi <= 8'h00;
		14'h259e:	ff_dbi <= 8'h00;
		14'h259f:	ff_dbi <= 8'h00;
		14'h25a0:	ff_dbi <= 8'h00;
		14'h25a1:	ff_dbi <= 8'h00;
		14'h25a2:	ff_dbi <= 8'h00;
		14'h25a3:	ff_dbi <= 8'h00;
		14'h25a4:	ff_dbi <= 8'h00;
		14'h25a5:	ff_dbi <= 8'h00;
		14'h25a6:	ff_dbi <= 8'h00;
		14'h25a7:	ff_dbi <= 8'h00;
		14'h25a8:	ff_dbi <= 8'h00;
		14'h25a9:	ff_dbi <= 8'h00;
		14'h25aa:	ff_dbi <= 8'h00;
		14'h25ab:	ff_dbi <= 8'h00;
		14'h25ac:	ff_dbi <= 8'h00;
		14'h25ad:	ff_dbi <= 8'h00;
		14'h25ae:	ff_dbi <= 8'h00;
		14'h25af:	ff_dbi <= 8'h00;
		14'h25b0:	ff_dbi <= 8'h00;
		14'h25b1:	ff_dbi <= 8'h00;
		14'h25b2:	ff_dbi <= 8'h00;
		14'h25b3:	ff_dbi <= 8'h00;
		14'h25b4:	ff_dbi <= 8'h00;
		14'h25b5:	ff_dbi <= 8'h00;
		14'h25b6:	ff_dbi <= 8'h00;
		14'h25b7:	ff_dbi <= 8'h00;
		14'h25b8:	ff_dbi <= 8'h00;
		14'h25b9:	ff_dbi <= 8'h00;
		14'h25ba:	ff_dbi <= 8'h00;
		14'h25bb:	ff_dbi <= 8'h00;
		14'h25bc:	ff_dbi <= 8'h00;
		14'h25bd:	ff_dbi <= 8'h00;
		14'h25be:	ff_dbi <= 8'h00;
		14'h25bf:	ff_dbi <= 8'h00;
		14'h25c0:	ff_dbi <= 8'h00;
		14'h25c1:	ff_dbi <= 8'h00;
		14'h25c2:	ff_dbi <= 8'h00;
		14'h25c3:	ff_dbi <= 8'h00;
		14'h25c4:	ff_dbi <= 8'h00;
		14'h25c5:	ff_dbi <= 8'h00;
		14'h25c6:	ff_dbi <= 8'h00;
		14'h25c7:	ff_dbi <= 8'h00;
		14'h25c8:	ff_dbi <= 8'h00;
		14'h25c9:	ff_dbi <= 8'h00;
		14'h25ca:	ff_dbi <= 8'h00;
		14'h25cb:	ff_dbi <= 8'h00;
		14'h25cc:	ff_dbi <= 8'h00;
		14'h25cd:	ff_dbi <= 8'h00;
		14'h25ce:	ff_dbi <= 8'h00;
		14'h25cf:	ff_dbi <= 8'h00;
		14'h25d0:	ff_dbi <= 8'h00;
		14'h25d1:	ff_dbi <= 8'h00;
		14'h25d2:	ff_dbi <= 8'h00;
		14'h25d3:	ff_dbi <= 8'h00;
		14'h25d4:	ff_dbi <= 8'h00;
		14'h25d5:	ff_dbi <= 8'h00;
		14'h25d6:	ff_dbi <= 8'h00;
		14'h25d7:	ff_dbi <= 8'h00;
		14'h25d8:	ff_dbi <= 8'h00;
		14'h25d9:	ff_dbi <= 8'h00;
		14'h25da:	ff_dbi <= 8'h00;
		14'h25db:	ff_dbi <= 8'h00;
		14'h25dc:	ff_dbi <= 8'h00;
		14'h25dd:	ff_dbi <= 8'h00;
		14'h25de:	ff_dbi <= 8'h00;
		14'h25df:	ff_dbi <= 8'h00;
		14'h25e0:	ff_dbi <= 8'h00;
		14'h25e1:	ff_dbi <= 8'h00;
		14'h25e2:	ff_dbi <= 8'h00;
		14'h25e3:	ff_dbi <= 8'h00;
		14'h25e4:	ff_dbi <= 8'h00;
		14'h25e5:	ff_dbi <= 8'h00;
		14'h25e6:	ff_dbi <= 8'h00;
		14'h25e7:	ff_dbi <= 8'h00;
		14'h25e8:	ff_dbi <= 8'h00;
		14'h25e9:	ff_dbi <= 8'h00;
		14'h25ea:	ff_dbi <= 8'h00;
		14'h25eb:	ff_dbi <= 8'h00;
		14'h25ec:	ff_dbi <= 8'h00;
		14'h25ed:	ff_dbi <= 8'h00;
		14'h25ee:	ff_dbi <= 8'h00;
		14'h25ef:	ff_dbi <= 8'h00;
		14'h25f0:	ff_dbi <= 8'h00;
		14'h25f1:	ff_dbi <= 8'h00;
		14'h25f2:	ff_dbi <= 8'h00;
		14'h25f3:	ff_dbi <= 8'h00;
		14'h25f4:	ff_dbi <= 8'h00;
		14'h25f5:	ff_dbi <= 8'h00;
		14'h25f6:	ff_dbi <= 8'h00;
		14'h25f7:	ff_dbi <= 8'h00;
		14'h25f8:	ff_dbi <= 8'h00;
		14'h25f9:	ff_dbi <= 8'h00;
		14'h25fa:	ff_dbi <= 8'h00;
		14'h25fb:	ff_dbi <= 8'h00;
		14'h25fc:	ff_dbi <= 8'h00;
		14'h25fd:	ff_dbi <= 8'h00;
		14'h25fe:	ff_dbi <= 8'h00;
		14'h25ff:	ff_dbi <= 8'h00;
		14'h2600:	ff_dbi <= 8'h00;
		14'h2601:	ff_dbi <= 8'h00;
		14'h2602:	ff_dbi <= 8'h00;
		14'h2603:	ff_dbi <= 8'h00;
		14'h2604:	ff_dbi <= 8'h00;
		14'h2605:	ff_dbi <= 8'h00;
		14'h2606:	ff_dbi <= 8'h00;
		14'h2607:	ff_dbi <= 8'h00;
		14'h2608:	ff_dbi <= 8'h00;
		14'h2609:	ff_dbi <= 8'h00;
		14'h260a:	ff_dbi <= 8'h00;
		14'h260b:	ff_dbi <= 8'h00;
		14'h260c:	ff_dbi <= 8'h00;
		14'h260d:	ff_dbi <= 8'h00;
		14'h260e:	ff_dbi <= 8'h00;
		14'h260f:	ff_dbi <= 8'h00;
		14'h2610:	ff_dbi <= 8'h00;
		14'h2611:	ff_dbi <= 8'h00;
		14'h2612:	ff_dbi <= 8'h00;
		14'h2613:	ff_dbi <= 8'h00;
		14'h2614:	ff_dbi <= 8'h00;
		14'h2615:	ff_dbi <= 8'h00;
		14'h2616:	ff_dbi <= 8'h00;
		14'h2617:	ff_dbi <= 8'h00;
		14'h2618:	ff_dbi <= 8'h00;
		14'h2619:	ff_dbi <= 8'h00;
		14'h261a:	ff_dbi <= 8'h00;
		14'h261b:	ff_dbi <= 8'h00;
		14'h261c:	ff_dbi <= 8'h00;
		14'h261d:	ff_dbi <= 8'h00;
		14'h261e:	ff_dbi <= 8'h00;
		14'h261f:	ff_dbi <= 8'h00;
		14'h2620:	ff_dbi <= 8'h00;
		14'h2621:	ff_dbi <= 8'h00;
		14'h2622:	ff_dbi <= 8'h00;
		14'h2623:	ff_dbi <= 8'h00;
		14'h2624:	ff_dbi <= 8'h00;
		14'h2625:	ff_dbi <= 8'h00;
		14'h2626:	ff_dbi <= 8'h00;
		14'h2627:	ff_dbi <= 8'h00;
		14'h2628:	ff_dbi <= 8'h00;
		14'h2629:	ff_dbi <= 8'h00;
		14'h262a:	ff_dbi <= 8'h00;
		14'h262b:	ff_dbi <= 8'h00;
		14'h262c:	ff_dbi <= 8'h00;
		14'h262d:	ff_dbi <= 8'h00;
		14'h262e:	ff_dbi <= 8'h00;
		14'h262f:	ff_dbi <= 8'h00;
		14'h2630:	ff_dbi <= 8'h00;
		14'h2631:	ff_dbi <= 8'h00;
		14'h2632:	ff_dbi <= 8'h00;
		14'h2633:	ff_dbi <= 8'h00;
		14'h2634:	ff_dbi <= 8'h00;
		14'h2635:	ff_dbi <= 8'h00;
		14'h2636:	ff_dbi <= 8'h00;
		14'h2637:	ff_dbi <= 8'h00;
		14'h2638:	ff_dbi <= 8'h00;
		14'h2639:	ff_dbi <= 8'h00;
		14'h263a:	ff_dbi <= 8'h00;
		14'h263b:	ff_dbi <= 8'h00;
		14'h263c:	ff_dbi <= 8'h00;
		14'h263d:	ff_dbi <= 8'h00;
		14'h263e:	ff_dbi <= 8'h00;
		14'h263f:	ff_dbi <= 8'h00;
		14'h2640:	ff_dbi <= 8'h00;
		14'h2641:	ff_dbi <= 8'h00;
		14'h2642:	ff_dbi <= 8'h00;
		14'h2643:	ff_dbi <= 8'h00;
		14'h2644:	ff_dbi <= 8'h00;
		14'h2645:	ff_dbi <= 8'h00;
		14'h2646:	ff_dbi <= 8'h00;
		14'h2647:	ff_dbi <= 8'h00;
		14'h2648:	ff_dbi <= 8'h00;
		14'h2649:	ff_dbi <= 8'h00;
		14'h264a:	ff_dbi <= 8'h00;
		14'h264b:	ff_dbi <= 8'h00;
		14'h264c:	ff_dbi <= 8'h00;
		14'h264d:	ff_dbi <= 8'h00;
		14'h264e:	ff_dbi <= 8'h00;
		14'h264f:	ff_dbi <= 8'h00;
		14'h2650:	ff_dbi <= 8'h00;
		14'h2651:	ff_dbi <= 8'h00;
		14'h2652:	ff_dbi <= 8'h00;
		14'h2653:	ff_dbi <= 8'h00;
		14'h2654:	ff_dbi <= 8'h00;
		14'h2655:	ff_dbi <= 8'h00;
		14'h2656:	ff_dbi <= 8'h00;
		14'h2657:	ff_dbi <= 8'h00;
		14'h2658:	ff_dbi <= 8'h00;
		14'h2659:	ff_dbi <= 8'h00;
		14'h265a:	ff_dbi <= 8'h00;
		14'h265b:	ff_dbi <= 8'h00;
		14'h265c:	ff_dbi <= 8'h00;
		14'h265d:	ff_dbi <= 8'h00;
		14'h265e:	ff_dbi <= 8'h00;
		14'h265f:	ff_dbi <= 8'h00;
		14'h2660:	ff_dbi <= 8'h00;
		14'h2661:	ff_dbi <= 8'h00;
		14'h2662:	ff_dbi <= 8'h00;
		14'h2663:	ff_dbi <= 8'h00;
		14'h2664:	ff_dbi <= 8'h00;
		14'h2665:	ff_dbi <= 8'h00;
		14'h2666:	ff_dbi <= 8'h00;
		14'h2667:	ff_dbi <= 8'h00;
		14'h2668:	ff_dbi <= 8'h00;
		14'h2669:	ff_dbi <= 8'h00;
		14'h266a:	ff_dbi <= 8'h00;
		14'h266b:	ff_dbi <= 8'h00;
		14'h266c:	ff_dbi <= 8'h00;
		14'h266d:	ff_dbi <= 8'h00;
		14'h266e:	ff_dbi <= 8'h00;
		14'h266f:	ff_dbi <= 8'h00;
		14'h2670:	ff_dbi <= 8'h00;
		14'h2671:	ff_dbi <= 8'h00;
		14'h2672:	ff_dbi <= 8'h00;
		14'h2673:	ff_dbi <= 8'h00;
		14'h2674:	ff_dbi <= 8'h00;
		14'h2675:	ff_dbi <= 8'h00;
		14'h2676:	ff_dbi <= 8'h00;
		14'h2677:	ff_dbi <= 8'h00;
		14'h2678:	ff_dbi <= 8'h00;
		14'h2679:	ff_dbi <= 8'h00;
		14'h267a:	ff_dbi <= 8'h00;
		14'h267b:	ff_dbi <= 8'h00;
		14'h267c:	ff_dbi <= 8'h00;
		14'h267d:	ff_dbi <= 8'h00;
		14'h267e:	ff_dbi <= 8'h00;
		14'h267f:	ff_dbi <= 8'h00;
		14'h2680:	ff_dbi <= 8'h00;
		14'h2681:	ff_dbi <= 8'h00;
		14'h2682:	ff_dbi <= 8'h00;
		14'h2683:	ff_dbi <= 8'h00;
		14'h2684:	ff_dbi <= 8'h00;
		14'h2685:	ff_dbi <= 8'h00;
		14'h2686:	ff_dbi <= 8'h00;
		14'h2687:	ff_dbi <= 8'h00;
		14'h2688:	ff_dbi <= 8'h00;
		14'h2689:	ff_dbi <= 8'h00;
		14'h268a:	ff_dbi <= 8'h00;
		14'h268b:	ff_dbi <= 8'h00;
		14'h268c:	ff_dbi <= 8'h00;
		14'h268d:	ff_dbi <= 8'h00;
		14'h268e:	ff_dbi <= 8'h00;
		14'h268f:	ff_dbi <= 8'h00;
		14'h2690:	ff_dbi <= 8'h00;
		14'h2691:	ff_dbi <= 8'h00;
		14'h2692:	ff_dbi <= 8'h00;
		14'h2693:	ff_dbi <= 8'h00;
		14'h2694:	ff_dbi <= 8'h00;
		14'h2695:	ff_dbi <= 8'h00;
		14'h2696:	ff_dbi <= 8'h00;
		14'h2697:	ff_dbi <= 8'h00;
		14'h2698:	ff_dbi <= 8'h00;
		14'h2699:	ff_dbi <= 8'h00;
		14'h269a:	ff_dbi <= 8'h00;
		14'h269b:	ff_dbi <= 8'h00;
		14'h269c:	ff_dbi <= 8'h00;
		14'h269d:	ff_dbi <= 8'h00;
		14'h269e:	ff_dbi <= 8'h00;
		14'h269f:	ff_dbi <= 8'h00;
		14'h26a0:	ff_dbi <= 8'h00;
		14'h26a1:	ff_dbi <= 8'h00;
		14'h26a2:	ff_dbi <= 8'h00;
		14'h26a3:	ff_dbi <= 8'h00;
		14'h26a4:	ff_dbi <= 8'h00;
		14'h26a5:	ff_dbi <= 8'h00;
		14'h26a6:	ff_dbi <= 8'h00;
		14'h26a7:	ff_dbi <= 8'h00;
		14'h26a8:	ff_dbi <= 8'h00;
		14'h26a9:	ff_dbi <= 8'h00;
		14'h26aa:	ff_dbi <= 8'h00;
		14'h26ab:	ff_dbi <= 8'h00;
		14'h26ac:	ff_dbi <= 8'h00;
		14'h26ad:	ff_dbi <= 8'h00;
		14'h26ae:	ff_dbi <= 8'h00;
		14'h26af:	ff_dbi <= 8'h00;
		14'h26b0:	ff_dbi <= 8'h00;
		14'h26b1:	ff_dbi <= 8'h00;
		14'h26b2:	ff_dbi <= 8'h00;
		14'h26b3:	ff_dbi <= 8'h00;
		14'h26b4:	ff_dbi <= 8'h00;
		14'h26b5:	ff_dbi <= 8'h00;
		14'h26b6:	ff_dbi <= 8'h00;
		14'h26b7:	ff_dbi <= 8'h00;
		14'h26b8:	ff_dbi <= 8'h00;
		14'h26b9:	ff_dbi <= 8'h00;
		14'h26ba:	ff_dbi <= 8'h00;
		14'h26bb:	ff_dbi <= 8'h00;
		14'h26bc:	ff_dbi <= 8'h00;
		14'h26bd:	ff_dbi <= 8'h00;
		14'h26be:	ff_dbi <= 8'h00;
		14'h26bf:	ff_dbi <= 8'h00;
		14'h26c0:	ff_dbi <= 8'h00;
		14'h26c1:	ff_dbi <= 8'h00;
		14'h26c2:	ff_dbi <= 8'h00;
		14'h26c3:	ff_dbi <= 8'h00;
		14'h26c4:	ff_dbi <= 8'h00;
		14'h26c5:	ff_dbi <= 8'h00;
		14'h26c6:	ff_dbi <= 8'h00;
		14'h26c7:	ff_dbi <= 8'h00;
		14'h26c8:	ff_dbi <= 8'h00;
		14'h26c9:	ff_dbi <= 8'h00;
		14'h26ca:	ff_dbi <= 8'h00;
		14'h26cb:	ff_dbi <= 8'h00;
		14'h26cc:	ff_dbi <= 8'h00;
		14'h26cd:	ff_dbi <= 8'h00;
		14'h26ce:	ff_dbi <= 8'h00;
		14'h26cf:	ff_dbi <= 8'h00;
		14'h26d0:	ff_dbi <= 8'h00;
		14'h26d1:	ff_dbi <= 8'h00;
		14'h26d2:	ff_dbi <= 8'h00;
		14'h26d3:	ff_dbi <= 8'h00;
		14'h26d4:	ff_dbi <= 8'h00;
		14'h26d5:	ff_dbi <= 8'h00;
		14'h26d6:	ff_dbi <= 8'h00;
		14'h26d7:	ff_dbi <= 8'h00;
		14'h26d8:	ff_dbi <= 8'h00;
		14'h26d9:	ff_dbi <= 8'h00;
		14'h26da:	ff_dbi <= 8'h00;
		14'h26db:	ff_dbi <= 8'h00;
		14'h26dc:	ff_dbi <= 8'h00;
		14'h26dd:	ff_dbi <= 8'h00;
		14'h26de:	ff_dbi <= 8'h00;
		14'h26df:	ff_dbi <= 8'h00;
		14'h26e0:	ff_dbi <= 8'h00;
		14'h26e1:	ff_dbi <= 8'h00;
		14'h26e2:	ff_dbi <= 8'h00;
		14'h26e3:	ff_dbi <= 8'h00;
		14'h26e4:	ff_dbi <= 8'h00;
		14'h26e5:	ff_dbi <= 8'h00;
		14'h26e6:	ff_dbi <= 8'h00;
		14'h26e7:	ff_dbi <= 8'h00;
		14'h26e8:	ff_dbi <= 8'h00;
		14'h26e9:	ff_dbi <= 8'h00;
		14'h26ea:	ff_dbi <= 8'h00;
		14'h26eb:	ff_dbi <= 8'h00;
		14'h26ec:	ff_dbi <= 8'h00;
		14'h26ed:	ff_dbi <= 8'h00;
		14'h26ee:	ff_dbi <= 8'h00;
		14'h26ef:	ff_dbi <= 8'h00;
		14'h26f0:	ff_dbi <= 8'h00;
		14'h26f1:	ff_dbi <= 8'h00;
		14'h26f2:	ff_dbi <= 8'h00;
		14'h26f3:	ff_dbi <= 8'h00;
		14'h26f4:	ff_dbi <= 8'h00;
		14'h26f5:	ff_dbi <= 8'h00;
		14'h26f6:	ff_dbi <= 8'h00;
		14'h26f7:	ff_dbi <= 8'h00;
		14'h26f8:	ff_dbi <= 8'h00;
		14'h26f9:	ff_dbi <= 8'h00;
		14'h26fa:	ff_dbi <= 8'h00;
		14'h26fb:	ff_dbi <= 8'h00;
		14'h26fc:	ff_dbi <= 8'h00;
		14'h26fd:	ff_dbi <= 8'h00;
		14'h26fe:	ff_dbi <= 8'h00;
		14'h26ff:	ff_dbi <= 8'h00;
		14'h2700:	ff_dbi <= 8'h00;
		14'h2701:	ff_dbi <= 8'h00;
		14'h2702:	ff_dbi <= 8'h00;
		14'h2703:	ff_dbi <= 8'h00;
		14'h2704:	ff_dbi <= 8'h00;
		14'h2705:	ff_dbi <= 8'h00;
		14'h2706:	ff_dbi <= 8'h00;
		14'h2707:	ff_dbi <= 8'h00;
		14'h2708:	ff_dbi <= 8'h00;
		14'h2709:	ff_dbi <= 8'h00;
		14'h270a:	ff_dbi <= 8'h00;
		14'h270b:	ff_dbi <= 8'h00;
		14'h270c:	ff_dbi <= 8'h00;
		14'h270d:	ff_dbi <= 8'h00;
		14'h270e:	ff_dbi <= 8'h00;
		14'h270f:	ff_dbi <= 8'h00;
		14'h2710:	ff_dbi <= 8'h00;
		14'h2711:	ff_dbi <= 8'h00;
		14'h2712:	ff_dbi <= 8'h00;
		14'h2713:	ff_dbi <= 8'h00;
		14'h2714:	ff_dbi <= 8'h00;
		14'h2715:	ff_dbi <= 8'h00;
		14'h2716:	ff_dbi <= 8'h00;
		14'h2717:	ff_dbi <= 8'h00;
		14'h2718:	ff_dbi <= 8'h00;
		14'h2719:	ff_dbi <= 8'h00;
		14'h271a:	ff_dbi <= 8'h00;
		14'h271b:	ff_dbi <= 8'h00;
		14'h271c:	ff_dbi <= 8'h00;
		14'h271d:	ff_dbi <= 8'h00;
		14'h271e:	ff_dbi <= 8'h00;
		14'h271f:	ff_dbi <= 8'h00;
		14'h2720:	ff_dbi <= 8'h00;
		14'h2721:	ff_dbi <= 8'h00;
		14'h2722:	ff_dbi <= 8'h00;
		14'h2723:	ff_dbi <= 8'h00;
		14'h2724:	ff_dbi <= 8'h00;
		14'h2725:	ff_dbi <= 8'h00;
		14'h2726:	ff_dbi <= 8'h00;
		14'h2727:	ff_dbi <= 8'h00;
		14'h2728:	ff_dbi <= 8'h00;
		14'h2729:	ff_dbi <= 8'h00;
		14'h272a:	ff_dbi <= 8'h00;
		14'h272b:	ff_dbi <= 8'h00;
		14'h272c:	ff_dbi <= 8'h00;
		14'h272d:	ff_dbi <= 8'h00;
		14'h272e:	ff_dbi <= 8'h00;
		14'h272f:	ff_dbi <= 8'h00;
		14'h2730:	ff_dbi <= 8'h00;
		14'h2731:	ff_dbi <= 8'h00;
		14'h2732:	ff_dbi <= 8'h00;
		14'h2733:	ff_dbi <= 8'h00;
		14'h2734:	ff_dbi <= 8'h00;
		14'h2735:	ff_dbi <= 8'h00;
		14'h2736:	ff_dbi <= 8'h00;
		14'h2737:	ff_dbi <= 8'h00;
		14'h2738:	ff_dbi <= 8'h00;
		14'h2739:	ff_dbi <= 8'h00;
		14'h273a:	ff_dbi <= 8'h00;
		14'h273b:	ff_dbi <= 8'h00;
		14'h273c:	ff_dbi <= 8'h00;
		14'h273d:	ff_dbi <= 8'h00;
		14'h273e:	ff_dbi <= 8'h00;
		14'h273f:	ff_dbi <= 8'h00;
		14'h2740:	ff_dbi <= 8'h00;
		14'h2741:	ff_dbi <= 8'h00;
		14'h2742:	ff_dbi <= 8'h00;
		14'h2743:	ff_dbi <= 8'h00;
		14'h2744:	ff_dbi <= 8'h00;
		14'h2745:	ff_dbi <= 8'h00;
		14'h2746:	ff_dbi <= 8'h00;
		14'h2747:	ff_dbi <= 8'h00;
		14'h2748:	ff_dbi <= 8'h00;
		14'h2749:	ff_dbi <= 8'h00;
		14'h274a:	ff_dbi <= 8'h00;
		14'h274b:	ff_dbi <= 8'h00;
		14'h274c:	ff_dbi <= 8'h00;
		14'h274d:	ff_dbi <= 8'h00;
		14'h274e:	ff_dbi <= 8'h00;
		14'h274f:	ff_dbi <= 8'h00;
		14'h2750:	ff_dbi <= 8'h00;
		14'h2751:	ff_dbi <= 8'h00;
		14'h2752:	ff_dbi <= 8'h00;
		14'h2753:	ff_dbi <= 8'h00;
		14'h2754:	ff_dbi <= 8'h00;
		14'h2755:	ff_dbi <= 8'h00;
		14'h2756:	ff_dbi <= 8'h00;
		14'h2757:	ff_dbi <= 8'h00;
		14'h2758:	ff_dbi <= 8'h00;
		14'h2759:	ff_dbi <= 8'h00;
		14'h275a:	ff_dbi <= 8'h00;
		14'h275b:	ff_dbi <= 8'h00;
		14'h275c:	ff_dbi <= 8'h00;
		14'h275d:	ff_dbi <= 8'h00;
		14'h275e:	ff_dbi <= 8'h00;
		14'h275f:	ff_dbi <= 8'h00;
		14'h2760:	ff_dbi <= 8'h00;
		14'h2761:	ff_dbi <= 8'h00;
		14'h2762:	ff_dbi <= 8'h00;
		14'h2763:	ff_dbi <= 8'h00;
		14'h2764:	ff_dbi <= 8'h00;
		14'h2765:	ff_dbi <= 8'h00;
		14'h2766:	ff_dbi <= 8'h00;
		14'h2767:	ff_dbi <= 8'h00;
		14'h2768:	ff_dbi <= 8'h00;
		14'h2769:	ff_dbi <= 8'h00;
		14'h276a:	ff_dbi <= 8'h00;
		14'h276b:	ff_dbi <= 8'h00;
		14'h276c:	ff_dbi <= 8'h00;
		14'h276d:	ff_dbi <= 8'h00;
		14'h276e:	ff_dbi <= 8'h00;
		14'h276f:	ff_dbi <= 8'h00;
		14'h2770:	ff_dbi <= 8'h00;
		14'h2771:	ff_dbi <= 8'h00;
		14'h2772:	ff_dbi <= 8'h00;
		14'h2773:	ff_dbi <= 8'h00;
		14'h2774:	ff_dbi <= 8'h00;
		14'h2775:	ff_dbi <= 8'h00;
		14'h2776:	ff_dbi <= 8'h00;
		14'h2777:	ff_dbi <= 8'h00;
		14'h2778:	ff_dbi <= 8'h00;
		14'h2779:	ff_dbi <= 8'h00;
		14'h277a:	ff_dbi <= 8'h00;
		14'h277b:	ff_dbi <= 8'h00;
		14'h277c:	ff_dbi <= 8'h00;
		14'h277d:	ff_dbi <= 8'h00;
		14'h277e:	ff_dbi <= 8'h00;
		14'h277f:	ff_dbi <= 8'h00;
		14'h2780:	ff_dbi <= 8'h00;
		14'h2781:	ff_dbi <= 8'h00;
		14'h2782:	ff_dbi <= 8'h00;
		14'h2783:	ff_dbi <= 8'h00;
		14'h2784:	ff_dbi <= 8'h00;
		14'h2785:	ff_dbi <= 8'h00;
		14'h2786:	ff_dbi <= 8'h00;
		14'h2787:	ff_dbi <= 8'h00;
		14'h2788:	ff_dbi <= 8'h00;
		14'h2789:	ff_dbi <= 8'h00;
		14'h278a:	ff_dbi <= 8'h00;
		14'h278b:	ff_dbi <= 8'h00;
		14'h278c:	ff_dbi <= 8'h00;
		14'h278d:	ff_dbi <= 8'h00;
		14'h278e:	ff_dbi <= 8'h00;
		14'h278f:	ff_dbi <= 8'h00;
		14'h2790:	ff_dbi <= 8'h00;
		14'h2791:	ff_dbi <= 8'h00;
		14'h2792:	ff_dbi <= 8'h00;
		14'h2793:	ff_dbi <= 8'h00;
		14'h2794:	ff_dbi <= 8'h00;
		14'h2795:	ff_dbi <= 8'h00;
		14'h2796:	ff_dbi <= 8'h00;
		14'h2797:	ff_dbi <= 8'h00;
		14'h2798:	ff_dbi <= 8'h00;
		14'h2799:	ff_dbi <= 8'h00;
		14'h279a:	ff_dbi <= 8'h00;
		14'h279b:	ff_dbi <= 8'h00;
		14'h279c:	ff_dbi <= 8'h00;
		14'h279d:	ff_dbi <= 8'h00;
		14'h279e:	ff_dbi <= 8'h00;
		14'h279f:	ff_dbi <= 8'h00;
		14'h27a0:	ff_dbi <= 8'h00;
		14'h27a1:	ff_dbi <= 8'h00;
		14'h27a2:	ff_dbi <= 8'h00;
		14'h27a3:	ff_dbi <= 8'h00;
		14'h27a4:	ff_dbi <= 8'h00;
		14'h27a5:	ff_dbi <= 8'h00;
		14'h27a6:	ff_dbi <= 8'h00;
		14'h27a7:	ff_dbi <= 8'h00;
		14'h27a8:	ff_dbi <= 8'h00;
		14'h27a9:	ff_dbi <= 8'h00;
		14'h27aa:	ff_dbi <= 8'h00;
		14'h27ab:	ff_dbi <= 8'h00;
		14'h27ac:	ff_dbi <= 8'h00;
		14'h27ad:	ff_dbi <= 8'h00;
		14'h27ae:	ff_dbi <= 8'h00;
		14'h27af:	ff_dbi <= 8'h00;
		14'h27b0:	ff_dbi <= 8'h00;
		14'h27b1:	ff_dbi <= 8'h00;
		14'h27b2:	ff_dbi <= 8'h00;
		14'h27b3:	ff_dbi <= 8'h00;
		14'h27b4:	ff_dbi <= 8'h00;
		14'h27b5:	ff_dbi <= 8'h00;
		14'h27b6:	ff_dbi <= 8'h00;
		14'h27b7:	ff_dbi <= 8'h00;
		14'h27b8:	ff_dbi <= 8'h00;
		14'h27b9:	ff_dbi <= 8'h00;
		14'h27ba:	ff_dbi <= 8'h00;
		14'h27bb:	ff_dbi <= 8'h00;
		14'h27bc:	ff_dbi <= 8'h00;
		14'h27bd:	ff_dbi <= 8'h00;
		14'h27be:	ff_dbi <= 8'h00;
		14'h27bf:	ff_dbi <= 8'h00;
		14'h27c0:	ff_dbi <= 8'h00;
		14'h27c1:	ff_dbi <= 8'h00;
		14'h27c2:	ff_dbi <= 8'h00;
		14'h27c3:	ff_dbi <= 8'h00;
		14'h27c4:	ff_dbi <= 8'h00;
		14'h27c5:	ff_dbi <= 8'h00;
		14'h27c6:	ff_dbi <= 8'h00;
		14'h27c7:	ff_dbi <= 8'h00;
		14'h27c8:	ff_dbi <= 8'h00;
		14'h27c9:	ff_dbi <= 8'h00;
		14'h27ca:	ff_dbi <= 8'h00;
		14'h27cb:	ff_dbi <= 8'h00;
		14'h27cc:	ff_dbi <= 8'h00;
		14'h27cd:	ff_dbi <= 8'h00;
		14'h27ce:	ff_dbi <= 8'h00;
		14'h27cf:	ff_dbi <= 8'h00;
		14'h27d0:	ff_dbi <= 8'h00;
		14'h27d1:	ff_dbi <= 8'h00;
		14'h27d2:	ff_dbi <= 8'h00;
		14'h27d3:	ff_dbi <= 8'h00;
		14'h27d4:	ff_dbi <= 8'h00;
		14'h27d5:	ff_dbi <= 8'h00;
		14'h27d6:	ff_dbi <= 8'h00;
		14'h27d7:	ff_dbi <= 8'h00;
		14'h27d8:	ff_dbi <= 8'h00;
		14'h27d9:	ff_dbi <= 8'h00;
		14'h27da:	ff_dbi <= 8'h00;
		14'h27db:	ff_dbi <= 8'h00;
		14'h27dc:	ff_dbi <= 8'h00;
		14'h27dd:	ff_dbi <= 8'h00;
		14'h27de:	ff_dbi <= 8'h00;
		14'h27df:	ff_dbi <= 8'h00;
		14'h27e0:	ff_dbi <= 8'h00;
		14'h27e1:	ff_dbi <= 8'h00;
		14'h27e2:	ff_dbi <= 8'h00;
		14'h27e3:	ff_dbi <= 8'h00;
		14'h27e4:	ff_dbi <= 8'h00;
		14'h27e5:	ff_dbi <= 8'h00;
		14'h27e6:	ff_dbi <= 8'h00;
		14'h27e7:	ff_dbi <= 8'h00;
		14'h27e8:	ff_dbi <= 8'h00;
		14'h27e9:	ff_dbi <= 8'h00;
		14'h27ea:	ff_dbi <= 8'h00;
		14'h27eb:	ff_dbi <= 8'h00;
		14'h27ec:	ff_dbi <= 8'h00;
		14'h27ed:	ff_dbi <= 8'h00;
		14'h27ee:	ff_dbi <= 8'h00;
		14'h27ef:	ff_dbi <= 8'h00;
		14'h27f0:	ff_dbi <= 8'h00;
		14'h27f1:	ff_dbi <= 8'h00;
		14'h27f2:	ff_dbi <= 8'h00;
		14'h27f3:	ff_dbi <= 8'h00;
		14'h27f4:	ff_dbi <= 8'h00;
		14'h27f5:	ff_dbi <= 8'h00;
		14'h27f6:	ff_dbi <= 8'h00;
		14'h27f7:	ff_dbi <= 8'h00;
		14'h27f8:	ff_dbi <= 8'h00;
		14'h27f9:	ff_dbi <= 8'h00;
		14'h27fa:	ff_dbi <= 8'h00;
		14'h27fb:	ff_dbi <= 8'h00;
		14'h27fc:	ff_dbi <= 8'h00;
		14'h27fd:	ff_dbi <= 8'h00;
		14'h27fe:	ff_dbi <= 8'h00;
		14'h27ff:	ff_dbi <= 8'h00;
		14'h2800:	ff_dbi <= 8'h00;
		14'h2801:	ff_dbi <= 8'h00;
		14'h2802:	ff_dbi <= 8'h00;
		14'h2803:	ff_dbi <= 8'h00;
		14'h2804:	ff_dbi <= 8'h00;
		14'h2805:	ff_dbi <= 8'h00;
		14'h2806:	ff_dbi <= 8'h00;
		14'h2807:	ff_dbi <= 8'h00;
		14'h2808:	ff_dbi <= 8'h00;
		14'h2809:	ff_dbi <= 8'h00;
		14'h280a:	ff_dbi <= 8'h00;
		14'h280b:	ff_dbi <= 8'h00;
		14'h280c:	ff_dbi <= 8'h00;
		14'h280d:	ff_dbi <= 8'h00;
		14'h280e:	ff_dbi <= 8'h00;
		14'h280f:	ff_dbi <= 8'h00;
		14'h2810:	ff_dbi <= 8'h00;
		14'h2811:	ff_dbi <= 8'h00;
		14'h2812:	ff_dbi <= 8'h00;
		14'h2813:	ff_dbi <= 8'h00;
		14'h2814:	ff_dbi <= 8'h00;
		14'h2815:	ff_dbi <= 8'h00;
		14'h2816:	ff_dbi <= 8'h00;
		14'h2817:	ff_dbi <= 8'h00;
		14'h2818:	ff_dbi <= 8'h00;
		14'h2819:	ff_dbi <= 8'h00;
		14'h281a:	ff_dbi <= 8'h00;
		14'h281b:	ff_dbi <= 8'h00;
		14'h281c:	ff_dbi <= 8'h00;
		14'h281d:	ff_dbi <= 8'h00;
		14'h281e:	ff_dbi <= 8'h00;
		14'h281f:	ff_dbi <= 8'h00;
		14'h2820:	ff_dbi <= 8'h00;
		14'h2821:	ff_dbi <= 8'h00;
		14'h2822:	ff_dbi <= 8'h00;
		14'h2823:	ff_dbi <= 8'h00;
		14'h2824:	ff_dbi <= 8'h00;
		14'h2825:	ff_dbi <= 8'h00;
		14'h2826:	ff_dbi <= 8'h00;
		14'h2827:	ff_dbi <= 8'h00;
		14'h2828:	ff_dbi <= 8'h00;
		14'h2829:	ff_dbi <= 8'h00;
		14'h282a:	ff_dbi <= 8'h00;
		14'h282b:	ff_dbi <= 8'h00;
		14'h282c:	ff_dbi <= 8'h00;
		14'h282d:	ff_dbi <= 8'h00;
		14'h282e:	ff_dbi <= 8'h00;
		14'h282f:	ff_dbi <= 8'h00;
		14'h2830:	ff_dbi <= 8'h00;
		14'h2831:	ff_dbi <= 8'h00;
		14'h2832:	ff_dbi <= 8'h00;
		14'h2833:	ff_dbi <= 8'h00;
		14'h2834:	ff_dbi <= 8'h00;
		14'h2835:	ff_dbi <= 8'h00;
		14'h2836:	ff_dbi <= 8'h00;
		14'h2837:	ff_dbi <= 8'h00;
		14'h2838:	ff_dbi <= 8'h00;
		14'h2839:	ff_dbi <= 8'h00;
		14'h283a:	ff_dbi <= 8'h00;
		14'h283b:	ff_dbi <= 8'h00;
		14'h283c:	ff_dbi <= 8'h00;
		14'h283d:	ff_dbi <= 8'h00;
		14'h283e:	ff_dbi <= 8'h00;
		14'h283f:	ff_dbi <= 8'h00;
		14'h2840:	ff_dbi <= 8'h00;
		14'h2841:	ff_dbi <= 8'h00;
		14'h2842:	ff_dbi <= 8'h00;
		14'h2843:	ff_dbi <= 8'h00;
		14'h2844:	ff_dbi <= 8'h00;
		14'h2845:	ff_dbi <= 8'h00;
		14'h2846:	ff_dbi <= 8'h00;
		14'h2847:	ff_dbi <= 8'h00;
		14'h2848:	ff_dbi <= 8'h00;
		14'h2849:	ff_dbi <= 8'h00;
		14'h284a:	ff_dbi <= 8'h00;
		14'h284b:	ff_dbi <= 8'h00;
		14'h284c:	ff_dbi <= 8'h00;
		14'h284d:	ff_dbi <= 8'h00;
		14'h284e:	ff_dbi <= 8'h00;
		14'h284f:	ff_dbi <= 8'h00;
		14'h2850:	ff_dbi <= 8'h00;
		14'h2851:	ff_dbi <= 8'h00;
		14'h2852:	ff_dbi <= 8'h00;
		14'h2853:	ff_dbi <= 8'h00;
		14'h2854:	ff_dbi <= 8'h00;
		14'h2855:	ff_dbi <= 8'h00;
		14'h2856:	ff_dbi <= 8'h00;
		14'h2857:	ff_dbi <= 8'h00;
		14'h2858:	ff_dbi <= 8'h00;
		14'h2859:	ff_dbi <= 8'h00;
		14'h285a:	ff_dbi <= 8'h00;
		14'h285b:	ff_dbi <= 8'h00;
		14'h285c:	ff_dbi <= 8'h00;
		14'h285d:	ff_dbi <= 8'h00;
		14'h285e:	ff_dbi <= 8'h00;
		14'h285f:	ff_dbi <= 8'h00;
		14'h2860:	ff_dbi <= 8'h00;
		14'h2861:	ff_dbi <= 8'h00;
		14'h2862:	ff_dbi <= 8'h00;
		14'h2863:	ff_dbi <= 8'h00;
		14'h2864:	ff_dbi <= 8'h00;
		14'h2865:	ff_dbi <= 8'h00;
		14'h2866:	ff_dbi <= 8'h00;
		14'h2867:	ff_dbi <= 8'h00;
		14'h2868:	ff_dbi <= 8'h00;
		14'h2869:	ff_dbi <= 8'h00;
		14'h286a:	ff_dbi <= 8'h00;
		14'h286b:	ff_dbi <= 8'h00;
		14'h286c:	ff_dbi <= 8'h00;
		14'h286d:	ff_dbi <= 8'h00;
		14'h286e:	ff_dbi <= 8'h00;
		14'h286f:	ff_dbi <= 8'h00;
		14'h2870:	ff_dbi <= 8'h00;
		14'h2871:	ff_dbi <= 8'h00;
		14'h2872:	ff_dbi <= 8'h00;
		14'h2873:	ff_dbi <= 8'h00;
		14'h2874:	ff_dbi <= 8'h00;
		14'h2875:	ff_dbi <= 8'h00;
		14'h2876:	ff_dbi <= 8'h00;
		14'h2877:	ff_dbi <= 8'h00;
		14'h2878:	ff_dbi <= 8'h00;
		14'h2879:	ff_dbi <= 8'h00;
		14'h287a:	ff_dbi <= 8'h00;
		14'h287b:	ff_dbi <= 8'h00;
		14'h287c:	ff_dbi <= 8'h00;
		14'h287d:	ff_dbi <= 8'h00;
		14'h287e:	ff_dbi <= 8'h00;
		14'h287f:	ff_dbi <= 8'h00;
		14'h2880:	ff_dbi <= 8'h00;
		14'h2881:	ff_dbi <= 8'h00;
		14'h2882:	ff_dbi <= 8'h00;
		14'h2883:	ff_dbi <= 8'h00;
		14'h2884:	ff_dbi <= 8'h00;
		14'h2885:	ff_dbi <= 8'h00;
		14'h2886:	ff_dbi <= 8'h00;
		14'h2887:	ff_dbi <= 8'h00;
		14'h2888:	ff_dbi <= 8'h00;
		14'h2889:	ff_dbi <= 8'h00;
		14'h288a:	ff_dbi <= 8'h00;
		14'h288b:	ff_dbi <= 8'h00;
		14'h288c:	ff_dbi <= 8'h00;
		14'h288d:	ff_dbi <= 8'h00;
		14'h288e:	ff_dbi <= 8'h00;
		14'h288f:	ff_dbi <= 8'h00;
		14'h2890:	ff_dbi <= 8'h00;
		14'h2891:	ff_dbi <= 8'h00;
		14'h2892:	ff_dbi <= 8'h00;
		14'h2893:	ff_dbi <= 8'h00;
		14'h2894:	ff_dbi <= 8'h00;
		14'h2895:	ff_dbi <= 8'h00;
		14'h2896:	ff_dbi <= 8'h00;
		14'h2897:	ff_dbi <= 8'h00;
		14'h2898:	ff_dbi <= 8'h00;
		14'h2899:	ff_dbi <= 8'h00;
		14'h289a:	ff_dbi <= 8'h00;
		14'h289b:	ff_dbi <= 8'h00;
		14'h289c:	ff_dbi <= 8'h00;
		14'h289d:	ff_dbi <= 8'h00;
		14'h289e:	ff_dbi <= 8'h00;
		14'h289f:	ff_dbi <= 8'h00;
		14'h28a0:	ff_dbi <= 8'h00;
		14'h28a1:	ff_dbi <= 8'h00;
		14'h28a2:	ff_dbi <= 8'h00;
		14'h28a3:	ff_dbi <= 8'h00;
		14'h28a4:	ff_dbi <= 8'h00;
		14'h28a5:	ff_dbi <= 8'h00;
		14'h28a6:	ff_dbi <= 8'h00;
		14'h28a7:	ff_dbi <= 8'h00;
		14'h28a8:	ff_dbi <= 8'h00;
		14'h28a9:	ff_dbi <= 8'h00;
		14'h28aa:	ff_dbi <= 8'h00;
		14'h28ab:	ff_dbi <= 8'h00;
		14'h28ac:	ff_dbi <= 8'h00;
		14'h28ad:	ff_dbi <= 8'h00;
		14'h28ae:	ff_dbi <= 8'h00;
		14'h28af:	ff_dbi <= 8'h00;
		14'h28b0:	ff_dbi <= 8'h00;
		14'h28b1:	ff_dbi <= 8'h00;
		14'h28b2:	ff_dbi <= 8'h00;
		14'h28b3:	ff_dbi <= 8'h00;
		14'h28b4:	ff_dbi <= 8'h00;
		14'h28b5:	ff_dbi <= 8'h00;
		14'h28b6:	ff_dbi <= 8'h00;
		14'h28b7:	ff_dbi <= 8'h00;
		14'h28b8:	ff_dbi <= 8'h00;
		14'h28b9:	ff_dbi <= 8'h00;
		14'h28ba:	ff_dbi <= 8'h00;
		14'h28bb:	ff_dbi <= 8'h00;
		14'h28bc:	ff_dbi <= 8'h00;
		14'h28bd:	ff_dbi <= 8'h00;
		14'h28be:	ff_dbi <= 8'h00;
		14'h28bf:	ff_dbi <= 8'h00;
		14'h28c0:	ff_dbi <= 8'h00;
		14'h28c1:	ff_dbi <= 8'h00;
		14'h28c2:	ff_dbi <= 8'h00;
		14'h28c3:	ff_dbi <= 8'h00;
		14'h28c4:	ff_dbi <= 8'h00;
		14'h28c5:	ff_dbi <= 8'h00;
		14'h28c6:	ff_dbi <= 8'h00;
		14'h28c7:	ff_dbi <= 8'h00;
		14'h28c8:	ff_dbi <= 8'h00;
		14'h28c9:	ff_dbi <= 8'h00;
		14'h28ca:	ff_dbi <= 8'h00;
		14'h28cb:	ff_dbi <= 8'h00;
		14'h28cc:	ff_dbi <= 8'h00;
		14'h28cd:	ff_dbi <= 8'h00;
		14'h28ce:	ff_dbi <= 8'h00;
		14'h28cf:	ff_dbi <= 8'h00;
		14'h28d0:	ff_dbi <= 8'h00;
		14'h28d1:	ff_dbi <= 8'h00;
		14'h28d2:	ff_dbi <= 8'h00;
		14'h28d3:	ff_dbi <= 8'h00;
		14'h28d4:	ff_dbi <= 8'h00;
		14'h28d5:	ff_dbi <= 8'h00;
		14'h28d6:	ff_dbi <= 8'h00;
		14'h28d7:	ff_dbi <= 8'h00;
		14'h28d8:	ff_dbi <= 8'h00;
		14'h28d9:	ff_dbi <= 8'h00;
		14'h28da:	ff_dbi <= 8'h00;
		14'h28db:	ff_dbi <= 8'h00;
		14'h28dc:	ff_dbi <= 8'h00;
		14'h28dd:	ff_dbi <= 8'h00;
		14'h28de:	ff_dbi <= 8'h00;
		14'h28df:	ff_dbi <= 8'h00;
		14'h28e0:	ff_dbi <= 8'h00;
		14'h28e1:	ff_dbi <= 8'h00;
		14'h28e2:	ff_dbi <= 8'h00;
		14'h28e3:	ff_dbi <= 8'h00;
		14'h28e4:	ff_dbi <= 8'h00;
		14'h28e5:	ff_dbi <= 8'h00;
		14'h28e6:	ff_dbi <= 8'h00;
		14'h28e7:	ff_dbi <= 8'h00;
		14'h28e8:	ff_dbi <= 8'h00;
		14'h28e9:	ff_dbi <= 8'h00;
		14'h28ea:	ff_dbi <= 8'h00;
		14'h28eb:	ff_dbi <= 8'h00;
		14'h28ec:	ff_dbi <= 8'h00;
		14'h28ed:	ff_dbi <= 8'h00;
		14'h28ee:	ff_dbi <= 8'h00;
		14'h28ef:	ff_dbi <= 8'h00;
		14'h28f0:	ff_dbi <= 8'h00;
		14'h28f1:	ff_dbi <= 8'h00;
		14'h28f2:	ff_dbi <= 8'h00;
		14'h28f3:	ff_dbi <= 8'h00;
		14'h28f4:	ff_dbi <= 8'h00;
		14'h28f5:	ff_dbi <= 8'h00;
		14'h28f6:	ff_dbi <= 8'h00;
		14'h28f7:	ff_dbi <= 8'h00;
		14'h28f8:	ff_dbi <= 8'h00;
		14'h28f9:	ff_dbi <= 8'h00;
		14'h28fa:	ff_dbi <= 8'h00;
		14'h28fb:	ff_dbi <= 8'h00;
		14'h28fc:	ff_dbi <= 8'h00;
		14'h28fd:	ff_dbi <= 8'h00;
		14'h28fe:	ff_dbi <= 8'h00;
		14'h28ff:	ff_dbi <= 8'h00;
		14'h2900:	ff_dbi <= 8'h00;
		14'h2901:	ff_dbi <= 8'h00;
		14'h2902:	ff_dbi <= 8'h00;
		14'h2903:	ff_dbi <= 8'h00;
		14'h2904:	ff_dbi <= 8'h00;
		14'h2905:	ff_dbi <= 8'h00;
		14'h2906:	ff_dbi <= 8'h00;
		14'h2907:	ff_dbi <= 8'h00;
		14'h2908:	ff_dbi <= 8'h00;
		14'h2909:	ff_dbi <= 8'h00;
		14'h290a:	ff_dbi <= 8'h00;
		14'h290b:	ff_dbi <= 8'h00;
		14'h290c:	ff_dbi <= 8'h00;
		14'h290d:	ff_dbi <= 8'h00;
		14'h290e:	ff_dbi <= 8'h00;
		14'h290f:	ff_dbi <= 8'h00;
		14'h2910:	ff_dbi <= 8'h00;
		14'h2911:	ff_dbi <= 8'h00;
		14'h2912:	ff_dbi <= 8'h00;
		14'h2913:	ff_dbi <= 8'h00;
		14'h2914:	ff_dbi <= 8'h00;
		14'h2915:	ff_dbi <= 8'h00;
		14'h2916:	ff_dbi <= 8'h00;
		14'h2917:	ff_dbi <= 8'h00;
		14'h2918:	ff_dbi <= 8'h00;
		14'h2919:	ff_dbi <= 8'h00;
		14'h291a:	ff_dbi <= 8'h00;
		14'h291b:	ff_dbi <= 8'h00;
		14'h291c:	ff_dbi <= 8'h00;
		14'h291d:	ff_dbi <= 8'h00;
		14'h291e:	ff_dbi <= 8'h00;
		14'h291f:	ff_dbi <= 8'h00;
		14'h2920:	ff_dbi <= 8'h00;
		14'h2921:	ff_dbi <= 8'h00;
		14'h2922:	ff_dbi <= 8'h00;
		14'h2923:	ff_dbi <= 8'h00;
		14'h2924:	ff_dbi <= 8'h00;
		14'h2925:	ff_dbi <= 8'h00;
		14'h2926:	ff_dbi <= 8'h00;
		14'h2927:	ff_dbi <= 8'h00;
		14'h2928:	ff_dbi <= 8'h00;
		14'h2929:	ff_dbi <= 8'h00;
		14'h292a:	ff_dbi <= 8'h00;
		14'h292b:	ff_dbi <= 8'h00;
		14'h292c:	ff_dbi <= 8'h00;
		14'h292d:	ff_dbi <= 8'h00;
		14'h292e:	ff_dbi <= 8'h00;
		14'h292f:	ff_dbi <= 8'h00;
		14'h2930:	ff_dbi <= 8'h00;
		14'h2931:	ff_dbi <= 8'h00;
		14'h2932:	ff_dbi <= 8'h00;
		14'h2933:	ff_dbi <= 8'h00;
		14'h2934:	ff_dbi <= 8'h00;
		14'h2935:	ff_dbi <= 8'h00;
		14'h2936:	ff_dbi <= 8'h00;
		14'h2937:	ff_dbi <= 8'h00;
		14'h2938:	ff_dbi <= 8'h00;
		14'h2939:	ff_dbi <= 8'h00;
		14'h293a:	ff_dbi <= 8'h00;
		14'h293b:	ff_dbi <= 8'h00;
		14'h293c:	ff_dbi <= 8'h00;
		14'h293d:	ff_dbi <= 8'h00;
		14'h293e:	ff_dbi <= 8'h00;
		14'h293f:	ff_dbi <= 8'h00;
		14'h2940:	ff_dbi <= 8'h00;
		14'h2941:	ff_dbi <= 8'h00;
		14'h2942:	ff_dbi <= 8'h00;
		14'h2943:	ff_dbi <= 8'h00;
		14'h2944:	ff_dbi <= 8'h00;
		14'h2945:	ff_dbi <= 8'h00;
		14'h2946:	ff_dbi <= 8'h00;
		14'h2947:	ff_dbi <= 8'h00;
		14'h2948:	ff_dbi <= 8'h00;
		14'h2949:	ff_dbi <= 8'h00;
		14'h294a:	ff_dbi <= 8'h00;
		14'h294b:	ff_dbi <= 8'h00;
		14'h294c:	ff_dbi <= 8'h00;
		14'h294d:	ff_dbi <= 8'h00;
		14'h294e:	ff_dbi <= 8'h00;
		14'h294f:	ff_dbi <= 8'h00;
		14'h2950:	ff_dbi <= 8'h00;
		14'h2951:	ff_dbi <= 8'h00;
		14'h2952:	ff_dbi <= 8'h00;
		14'h2953:	ff_dbi <= 8'h00;
		14'h2954:	ff_dbi <= 8'h00;
		14'h2955:	ff_dbi <= 8'h00;
		14'h2956:	ff_dbi <= 8'h00;
		14'h2957:	ff_dbi <= 8'h00;
		14'h2958:	ff_dbi <= 8'h00;
		14'h2959:	ff_dbi <= 8'h00;
		14'h295a:	ff_dbi <= 8'h00;
		14'h295b:	ff_dbi <= 8'h00;
		14'h295c:	ff_dbi <= 8'h00;
		14'h295d:	ff_dbi <= 8'h00;
		14'h295e:	ff_dbi <= 8'h00;
		14'h295f:	ff_dbi <= 8'h00;
		14'h2960:	ff_dbi <= 8'h00;
		14'h2961:	ff_dbi <= 8'h00;
		14'h2962:	ff_dbi <= 8'h00;
		14'h2963:	ff_dbi <= 8'h00;
		14'h2964:	ff_dbi <= 8'h00;
		14'h2965:	ff_dbi <= 8'h00;
		14'h2966:	ff_dbi <= 8'h00;
		14'h2967:	ff_dbi <= 8'h00;
		14'h2968:	ff_dbi <= 8'h00;
		14'h2969:	ff_dbi <= 8'h00;
		14'h296a:	ff_dbi <= 8'h00;
		14'h296b:	ff_dbi <= 8'h00;
		14'h296c:	ff_dbi <= 8'h00;
		14'h296d:	ff_dbi <= 8'h00;
		14'h296e:	ff_dbi <= 8'h00;
		14'h296f:	ff_dbi <= 8'h00;
		14'h2970:	ff_dbi <= 8'h00;
		14'h2971:	ff_dbi <= 8'h00;
		14'h2972:	ff_dbi <= 8'h00;
		14'h2973:	ff_dbi <= 8'h00;
		14'h2974:	ff_dbi <= 8'h00;
		14'h2975:	ff_dbi <= 8'h00;
		14'h2976:	ff_dbi <= 8'h00;
		14'h2977:	ff_dbi <= 8'h00;
		14'h2978:	ff_dbi <= 8'h00;
		14'h2979:	ff_dbi <= 8'h00;
		14'h297a:	ff_dbi <= 8'h00;
		14'h297b:	ff_dbi <= 8'h00;
		14'h297c:	ff_dbi <= 8'h00;
		14'h297d:	ff_dbi <= 8'h00;
		14'h297e:	ff_dbi <= 8'h00;
		14'h297f:	ff_dbi <= 8'h00;
		14'h2980:	ff_dbi <= 8'h00;
		14'h2981:	ff_dbi <= 8'h00;
		14'h2982:	ff_dbi <= 8'h00;
		14'h2983:	ff_dbi <= 8'h00;
		14'h2984:	ff_dbi <= 8'h00;
		14'h2985:	ff_dbi <= 8'h00;
		14'h2986:	ff_dbi <= 8'h00;
		14'h2987:	ff_dbi <= 8'h00;
		14'h2988:	ff_dbi <= 8'h00;
		14'h2989:	ff_dbi <= 8'h00;
		14'h298a:	ff_dbi <= 8'h00;
		14'h298b:	ff_dbi <= 8'h00;
		14'h298c:	ff_dbi <= 8'h00;
		14'h298d:	ff_dbi <= 8'h00;
		14'h298e:	ff_dbi <= 8'h00;
		14'h298f:	ff_dbi <= 8'h00;
		14'h2990:	ff_dbi <= 8'h00;
		14'h2991:	ff_dbi <= 8'h00;
		14'h2992:	ff_dbi <= 8'h00;
		14'h2993:	ff_dbi <= 8'h00;
		14'h2994:	ff_dbi <= 8'h00;
		14'h2995:	ff_dbi <= 8'h00;
		14'h2996:	ff_dbi <= 8'h00;
		14'h2997:	ff_dbi <= 8'h00;
		14'h2998:	ff_dbi <= 8'h00;
		14'h2999:	ff_dbi <= 8'h00;
		14'h299a:	ff_dbi <= 8'h00;
		14'h299b:	ff_dbi <= 8'h00;
		14'h299c:	ff_dbi <= 8'h00;
		14'h299d:	ff_dbi <= 8'h00;
		14'h299e:	ff_dbi <= 8'h00;
		14'h299f:	ff_dbi <= 8'h00;
		14'h29a0:	ff_dbi <= 8'h00;
		14'h29a1:	ff_dbi <= 8'h00;
		14'h29a2:	ff_dbi <= 8'h00;
		14'h29a3:	ff_dbi <= 8'h00;
		14'h29a4:	ff_dbi <= 8'h00;
		14'h29a5:	ff_dbi <= 8'h00;
		14'h29a6:	ff_dbi <= 8'h00;
		14'h29a7:	ff_dbi <= 8'h00;
		14'h29a8:	ff_dbi <= 8'h00;
		14'h29a9:	ff_dbi <= 8'h00;
		14'h29aa:	ff_dbi <= 8'h00;
		14'h29ab:	ff_dbi <= 8'h00;
		14'h29ac:	ff_dbi <= 8'h00;
		14'h29ad:	ff_dbi <= 8'h00;
		14'h29ae:	ff_dbi <= 8'h00;
		14'h29af:	ff_dbi <= 8'h00;
		14'h29b0:	ff_dbi <= 8'h00;
		14'h29b1:	ff_dbi <= 8'h00;
		14'h29b2:	ff_dbi <= 8'h00;
		14'h29b3:	ff_dbi <= 8'h00;
		14'h29b4:	ff_dbi <= 8'h00;
		14'h29b5:	ff_dbi <= 8'h00;
		14'h29b6:	ff_dbi <= 8'h00;
		14'h29b7:	ff_dbi <= 8'h00;
		14'h29b8:	ff_dbi <= 8'h00;
		14'h29b9:	ff_dbi <= 8'h00;
		14'h29ba:	ff_dbi <= 8'h00;
		14'h29bb:	ff_dbi <= 8'h00;
		14'h29bc:	ff_dbi <= 8'h00;
		14'h29bd:	ff_dbi <= 8'h00;
		14'h29be:	ff_dbi <= 8'h00;
		14'h29bf:	ff_dbi <= 8'h00;
		14'h29c0:	ff_dbi <= 8'h00;
		14'h29c1:	ff_dbi <= 8'h00;
		14'h29c2:	ff_dbi <= 8'h00;
		14'h29c3:	ff_dbi <= 8'h00;
		14'h29c4:	ff_dbi <= 8'h00;
		14'h29c5:	ff_dbi <= 8'h00;
		14'h29c6:	ff_dbi <= 8'h00;
		14'h29c7:	ff_dbi <= 8'h00;
		14'h29c8:	ff_dbi <= 8'h00;
		14'h29c9:	ff_dbi <= 8'h00;
		14'h29ca:	ff_dbi <= 8'h00;
		14'h29cb:	ff_dbi <= 8'h00;
		14'h29cc:	ff_dbi <= 8'h00;
		14'h29cd:	ff_dbi <= 8'h00;
		14'h29ce:	ff_dbi <= 8'h00;
		14'h29cf:	ff_dbi <= 8'h00;
		14'h29d0:	ff_dbi <= 8'h00;
		14'h29d1:	ff_dbi <= 8'h00;
		14'h29d2:	ff_dbi <= 8'h00;
		14'h29d3:	ff_dbi <= 8'h00;
		14'h29d4:	ff_dbi <= 8'h00;
		14'h29d5:	ff_dbi <= 8'h00;
		14'h29d6:	ff_dbi <= 8'h00;
		14'h29d7:	ff_dbi <= 8'h00;
		14'h29d8:	ff_dbi <= 8'h00;
		14'h29d9:	ff_dbi <= 8'h00;
		14'h29da:	ff_dbi <= 8'h00;
		14'h29db:	ff_dbi <= 8'h00;
		14'h29dc:	ff_dbi <= 8'h00;
		14'h29dd:	ff_dbi <= 8'h00;
		14'h29de:	ff_dbi <= 8'h00;
		14'h29df:	ff_dbi <= 8'h00;
		14'h29e0:	ff_dbi <= 8'h00;
		14'h29e1:	ff_dbi <= 8'h00;
		14'h29e2:	ff_dbi <= 8'h00;
		14'h29e3:	ff_dbi <= 8'h00;
		14'h29e4:	ff_dbi <= 8'h00;
		14'h29e5:	ff_dbi <= 8'h00;
		14'h29e6:	ff_dbi <= 8'h00;
		14'h29e7:	ff_dbi <= 8'h00;
		14'h29e8:	ff_dbi <= 8'h00;
		14'h29e9:	ff_dbi <= 8'h00;
		14'h29ea:	ff_dbi <= 8'h00;
		14'h29eb:	ff_dbi <= 8'h00;
		14'h29ec:	ff_dbi <= 8'h00;
		14'h29ed:	ff_dbi <= 8'h00;
		14'h29ee:	ff_dbi <= 8'h00;
		14'h29ef:	ff_dbi <= 8'h00;
		14'h29f0:	ff_dbi <= 8'h00;
		14'h29f1:	ff_dbi <= 8'h00;
		14'h29f2:	ff_dbi <= 8'h00;
		14'h29f3:	ff_dbi <= 8'h00;
		14'h29f4:	ff_dbi <= 8'h00;
		14'h29f5:	ff_dbi <= 8'h00;
		14'h29f6:	ff_dbi <= 8'h00;
		14'h29f7:	ff_dbi <= 8'h00;
		14'h29f8:	ff_dbi <= 8'h00;
		14'h29f9:	ff_dbi <= 8'h00;
		14'h29fa:	ff_dbi <= 8'h00;
		14'h29fb:	ff_dbi <= 8'h00;
		14'h29fc:	ff_dbi <= 8'h00;
		14'h29fd:	ff_dbi <= 8'h00;
		14'h29fe:	ff_dbi <= 8'h00;
		14'h29ff:	ff_dbi <= 8'h00;
		14'h2a00:	ff_dbi <= 8'h00;
		14'h2a01:	ff_dbi <= 8'h00;
		14'h2a02:	ff_dbi <= 8'h00;
		14'h2a03:	ff_dbi <= 8'h00;
		14'h2a04:	ff_dbi <= 8'h00;
		14'h2a05:	ff_dbi <= 8'h00;
		14'h2a06:	ff_dbi <= 8'h00;
		14'h2a07:	ff_dbi <= 8'h00;
		14'h2a08:	ff_dbi <= 8'h00;
		14'h2a09:	ff_dbi <= 8'h00;
		14'h2a0a:	ff_dbi <= 8'h00;
		14'h2a0b:	ff_dbi <= 8'h00;
		14'h2a0c:	ff_dbi <= 8'h00;
		14'h2a0d:	ff_dbi <= 8'h00;
		14'h2a0e:	ff_dbi <= 8'h00;
		14'h2a0f:	ff_dbi <= 8'h00;
		14'h2a10:	ff_dbi <= 8'h00;
		14'h2a11:	ff_dbi <= 8'h00;
		14'h2a12:	ff_dbi <= 8'h00;
		14'h2a13:	ff_dbi <= 8'h00;
		14'h2a14:	ff_dbi <= 8'h00;
		14'h2a15:	ff_dbi <= 8'h00;
		14'h2a16:	ff_dbi <= 8'h00;
		14'h2a17:	ff_dbi <= 8'h00;
		14'h2a18:	ff_dbi <= 8'h00;
		14'h2a19:	ff_dbi <= 8'h00;
		14'h2a1a:	ff_dbi <= 8'h00;
		14'h2a1b:	ff_dbi <= 8'h00;
		14'h2a1c:	ff_dbi <= 8'h00;
		14'h2a1d:	ff_dbi <= 8'h00;
		14'h2a1e:	ff_dbi <= 8'h00;
		14'h2a1f:	ff_dbi <= 8'h00;
		14'h2a20:	ff_dbi <= 8'h00;
		14'h2a21:	ff_dbi <= 8'h00;
		14'h2a22:	ff_dbi <= 8'h00;
		14'h2a23:	ff_dbi <= 8'h00;
		14'h2a24:	ff_dbi <= 8'h00;
		14'h2a25:	ff_dbi <= 8'h00;
		14'h2a26:	ff_dbi <= 8'h00;
		14'h2a27:	ff_dbi <= 8'h00;
		14'h2a28:	ff_dbi <= 8'h00;
		14'h2a29:	ff_dbi <= 8'h00;
		14'h2a2a:	ff_dbi <= 8'h00;
		14'h2a2b:	ff_dbi <= 8'h00;
		14'h2a2c:	ff_dbi <= 8'h00;
		14'h2a2d:	ff_dbi <= 8'h00;
		14'h2a2e:	ff_dbi <= 8'h00;
		14'h2a2f:	ff_dbi <= 8'h00;
		14'h2a30:	ff_dbi <= 8'h00;
		14'h2a31:	ff_dbi <= 8'h00;
		14'h2a32:	ff_dbi <= 8'h00;
		14'h2a33:	ff_dbi <= 8'h00;
		14'h2a34:	ff_dbi <= 8'h00;
		14'h2a35:	ff_dbi <= 8'h00;
		14'h2a36:	ff_dbi <= 8'h00;
		14'h2a37:	ff_dbi <= 8'h00;
		14'h2a38:	ff_dbi <= 8'h00;
		14'h2a39:	ff_dbi <= 8'h00;
		14'h2a3a:	ff_dbi <= 8'h00;
		14'h2a3b:	ff_dbi <= 8'h00;
		14'h2a3c:	ff_dbi <= 8'h00;
		14'h2a3d:	ff_dbi <= 8'h00;
		14'h2a3e:	ff_dbi <= 8'h00;
		14'h2a3f:	ff_dbi <= 8'h00;
		14'h2a40:	ff_dbi <= 8'h00;
		14'h2a41:	ff_dbi <= 8'h00;
		14'h2a42:	ff_dbi <= 8'h00;
		14'h2a43:	ff_dbi <= 8'h00;
		14'h2a44:	ff_dbi <= 8'h00;
		14'h2a45:	ff_dbi <= 8'h00;
		14'h2a46:	ff_dbi <= 8'h00;
		14'h2a47:	ff_dbi <= 8'h00;
		14'h2a48:	ff_dbi <= 8'h00;
		14'h2a49:	ff_dbi <= 8'h00;
		14'h2a4a:	ff_dbi <= 8'h00;
		14'h2a4b:	ff_dbi <= 8'h00;
		14'h2a4c:	ff_dbi <= 8'h00;
		14'h2a4d:	ff_dbi <= 8'h00;
		14'h2a4e:	ff_dbi <= 8'h00;
		14'h2a4f:	ff_dbi <= 8'h00;
		14'h2a50:	ff_dbi <= 8'h00;
		14'h2a51:	ff_dbi <= 8'h00;
		14'h2a52:	ff_dbi <= 8'h00;
		14'h2a53:	ff_dbi <= 8'h00;
		14'h2a54:	ff_dbi <= 8'h00;
		14'h2a55:	ff_dbi <= 8'h00;
		14'h2a56:	ff_dbi <= 8'h00;
		14'h2a57:	ff_dbi <= 8'h00;
		14'h2a58:	ff_dbi <= 8'h00;
		14'h2a59:	ff_dbi <= 8'h00;
		14'h2a5a:	ff_dbi <= 8'h00;
		14'h2a5b:	ff_dbi <= 8'h00;
		14'h2a5c:	ff_dbi <= 8'h00;
		14'h2a5d:	ff_dbi <= 8'h00;
		14'h2a5e:	ff_dbi <= 8'h00;
		14'h2a5f:	ff_dbi <= 8'h00;
		14'h2a60:	ff_dbi <= 8'h00;
		14'h2a61:	ff_dbi <= 8'h00;
		14'h2a62:	ff_dbi <= 8'h00;
		14'h2a63:	ff_dbi <= 8'h00;
		14'h2a64:	ff_dbi <= 8'h00;
		14'h2a65:	ff_dbi <= 8'h00;
		14'h2a66:	ff_dbi <= 8'h00;
		14'h2a67:	ff_dbi <= 8'h00;
		14'h2a68:	ff_dbi <= 8'h00;
		14'h2a69:	ff_dbi <= 8'h00;
		14'h2a6a:	ff_dbi <= 8'h00;
		14'h2a6b:	ff_dbi <= 8'h00;
		14'h2a6c:	ff_dbi <= 8'h00;
		14'h2a6d:	ff_dbi <= 8'h00;
		14'h2a6e:	ff_dbi <= 8'h00;
		14'h2a6f:	ff_dbi <= 8'h00;
		14'h2a70:	ff_dbi <= 8'h00;
		14'h2a71:	ff_dbi <= 8'h00;
		14'h2a72:	ff_dbi <= 8'h00;
		14'h2a73:	ff_dbi <= 8'h00;
		14'h2a74:	ff_dbi <= 8'h00;
		14'h2a75:	ff_dbi <= 8'h00;
		14'h2a76:	ff_dbi <= 8'h00;
		14'h2a77:	ff_dbi <= 8'h00;
		14'h2a78:	ff_dbi <= 8'h00;
		14'h2a79:	ff_dbi <= 8'h00;
		14'h2a7a:	ff_dbi <= 8'h00;
		14'h2a7b:	ff_dbi <= 8'h00;
		14'h2a7c:	ff_dbi <= 8'h00;
		14'h2a7d:	ff_dbi <= 8'h00;
		14'h2a7e:	ff_dbi <= 8'h00;
		14'h2a7f:	ff_dbi <= 8'h00;
		14'h2a80:	ff_dbi <= 8'h00;
		14'h2a81:	ff_dbi <= 8'h00;
		14'h2a82:	ff_dbi <= 8'h00;
		14'h2a83:	ff_dbi <= 8'h00;
		14'h2a84:	ff_dbi <= 8'h00;
		14'h2a85:	ff_dbi <= 8'h00;
		14'h2a86:	ff_dbi <= 8'h00;
		14'h2a87:	ff_dbi <= 8'h00;
		14'h2a88:	ff_dbi <= 8'h00;
		14'h2a89:	ff_dbi <= 8'h00;
		14'h2a8a:	ff_dbi <= 8'h00;
		14'h2a8b:	ff_dbi <= 8'h00;
		14'h2a8c:	ff_dbi <= 8'h00;
		14'h2a8d:	ff_dbi <= 8'h00;
		14'h2a8e:	ff_dbi <= 8'h00;
		14'h2a8f:	ff_dbi <= 8'h00;
		14'h2a90:	ff_dbi <= 8'h00;
		14'h2a91:	ff_dbi <= 8'h00;
		14'h2a92:	ff_dbi <= 8'h00;
		14'h2a93:	ff_dbi <= 8'h00;
		14'h2a94:	ff_dbi <= 8'h00;
		14'h2a95:	ff_dbi <= 8'h00;
		14'h2a96:	ff_dbi <= 8'h00;
		14'h2a97:	ff_dbi <= 8'h00;
		14'h2a98:	ff_dbi <= 8'h00;
		14'h2a99:	ff_dbi <= 8'h00;
		14'h2a9a:	ff_dbi <= 8'h00;
		14'h2a9b:	ff_dbi <= 8'h00;
		14'h2a9c:	ff_dbi <= 8'h00;
		14'h2a9d:	ff_dbi <= 8'h00;
		14'h2a9e:	ff_dbi <= 8'h00;
		14'h2a9f:	ff_dbi <= 8'h00;
		14'h2aa0:	ff_dbi <= 8'h00;
		14'h2aa1:	ff_dbi <= 8'h00;
		14'h2aa2:	ff_dbi <= 8'h00;
		14'h2aa3:	ff_dbi <= 8'h00;
		14'h2aa4:	ff_dbi <= 8'h00;
		14'h2aa5:	ff_dbi <= 8'h00;
		14'h2aa6:	ff_dbi <= 8'h00;
		14'h2aa7:	ff_dbi <= 8'h00;
		14'h2aa8:	ff_dbi <= 8'h00;
		14'h2aa9:	ff_dbi <= 8'h00;
		14'h2aaa:	ff_dbi <= 8'h00;
		14'h2aab:	ff_dbi <= 8'h00;
		14'h2aac:	ff_dbi <= 8'h00;
		14'h2aad:	ff_dbi <= 8'h00;
		14'h2aae:	ff_dbi <= 8'h00;
		14'h2aaf:	ff_dbi <= 8'h00;
		14'h2ab0:	ff_dbi <= 8'h00;
		14'h2ab1:	ff_dbi <= 8'h00;
		14'h2ab2:	ff_dbi <= 8'h00;
		14'h2ab3:	ff_dbi <= 8'h00;
		14'h2ab4:	ff_dbi <= 8'h00;
		14'h2ab5:	ff_dbi <= 8'h00;
		14'h2ab6:	ff_dbi <= 8'h00;
		14'h2ab7:	ff_dbi <= 8'h00;
		14'h2ab8:	ff_dbi <= 8'h00;
		14'h2ab9:	ff_dbi <= 8'h00;
		14'h2aba:	ff_dbi <= 8'h00;
		14'h2abb:	ff_dbi <= 8'h00;
		14'h2abc:	ff_dbi <= 8'h00;
		14'h2abd:	ff_dbi <= 8'h00;
		14'h2abe:	ff_dbi <= 8'h00;
		14'h2abf:	ff_dbi <= 8'h00;
		14'h2ac0:	ff_dbi <= 8'h00;
		14'h2ac1:	ff_dbi <= 8'h00;
		14'h2ac2:	ff_dbi <= 8'h00;
		14'h2ac3:	ff_dbi <= 8'h00;
		14'h2ac4:	ff_dbi <= 8'h00;
		14'h2ac5:	ff_dbi <= 8'h00;
		14'h2ac6:	ff_dbi <= 8'h00;
		14'h2ac7:	ff_dbi <= 8'h00;
		14'h2ac8:	ff_dbi <= 8'h00;
		14'h2ac9:	ff_dbi <= 8'h00;
		14'h2aca:	ff_dbi <= 8'h00;
		14'h2acb:	ff_dbi <= 8'h00;
		14'h2acc:	ff_dbi <= 8'h00;
		14'h2acd:	ff_dbi <= 8'h00;
		14'h2ace:	ff_dbi <= 8'h00;
		14'h2acf:	ff_dbi <= 8'h00;
		14'h2ad0:	ff_dbi <= 8'h00;
		14'h2ad1:	ff_dbi <= 8'h00;
		14'h2ad2:	ff_dbi <= 8'h00;
		14'h2ad3:	ff_dbi <= 8'h00;
		14'h2ad4:	ff_dbi <= 8'h00;
		14'h2ad5:	ff_dbi <= 8'h00;
		14'h2ad6:	ff_dbi <= 8'h00;
		14'h2ad7:	ff_dbi <= 8'h00;
		14'h2ad8:	ff_dbi <= 8'h00;
		14'h2ad9:	ff_dbi <= 8'h00;
		14'h2ada:	ff_dbi <= 8'h00;
		14'h2adb:	ff_dbi <= 8'h00;
		14'h2adc:	ff_dbi <= 8'h00;
		14'h2add:	ff_dbi <= 8'h00;
		14'h2ade:	ff_dbi <= 8'h00;
		14'h2adf:	ff_dbi <= 8'h00;
		14'h2ae0:	ff_dbi <= 8'h00;
		14'h2ae1:	ff_dbi <= 8'h00;
		14'h2ae2:	ff_dbi <= 8'h00;
		14'h2ae3:	ff_dbi <= 8'h00;
		14'h2ae4:	ff_dbi <= 8'h00;
		14'h2ae5:	ff_dbi <= 8'h00;
		14'h2ae6:	ff_dbi <= 8'h00;
		14'h2ae7:	ff_dbi <= 8'h00;
		14'h2ae8:	ff_dbi <= 8'h00;
		14'h2ae9:	ff_dbi <= 8'h00;
		14'h2aea:	ff_dbi <= 8'h00;
		14'h2aeb:	ff_dbi <= 8'h00;
		14'h2aec:	ff_dbi <= 8'h00;
		14'h2aed:	ff_dbi <= 8'h00;
		14'h2aee:	ff_dbi <= 8'h00;
		14'h2aef:	ff_dbi <= 8'h00;
		14'h2af0:	ff_dbi <= 8'h00;
		14'h2af1:	ff_dbi <= 8'h00;
		14'h2af2:	ff_dbi <= 8'h00;
		14'h2af3:	ff_dbi <= 8'h00;
		14'h2af4:	ff_dbi <= 8'h00;
		14'h2af5:	ff_dbi <= 8'h00;
		14'h2af6:	ff_dbi <= 8'h00;
		14'h2af7:	ff_dbi <= 8'h00;
		14'h2af8:	ff_dbi <= 8'h00;
		14'h2af9:	ff_dbi <= 8'h00;
		14'h2afa:	ff_dbi <= 8'h00;
		14'h2afb:	ff_dbi <= 8'h00;
		14'h2afc:	ff_dbi <= 8'h00;
		14'h2afd:	ff_dbi <= 8'h00;
		14'h2afe:	ff_dbi <= 8'h00;
		14'h2aff:	ff_dbi <= 8'h00;
		14'h2b00:	ff_dbi <= 8'h00;
		14'h2b01:	ff_dbi <= 8'h00;
		14'h2b02:	ff_dbi <= 8'h00;
		14'h2b03:	ff_dbi <= 8'h00;
		14'h2b04:	ff_dbi <= 8'h00;
		14'h2b05:	ff_dbi <= 8'h00;
		14'h2b06:	ff_dbi <= 8'h00;
		14'h2b07:	ff_dbi <= 8'h00;
		14'h2b08:	ff_dbi <= 8'h00;
		14'h2b09:	ff_dbi <= 8'h00;
		14'h2b0a:	ff_dbi <= 8'h00;
		14'h2b0b:	ff_dbi <= 8'h00;
		14'h2b0c:	ff_dbi <= 8'h00;
		14'h2b0d:	ff_dbi <= 8'h00;
		14'h2b0e:	ff_dbi <= 8'h00;
		14'h2b0f:	ff_dbi <= 8'h00;
		14'h2b10:	ff_dbi <= 8'h00;
		14'h2b11:	ff_dbi <= 8'h00;
		14'h2b12:	ff_dbi <= 8'h00;
		14'h2b13:	ff_dbi <= 8'h00;
		14'h2b14:	ff_dbi <= 8'h00;
		14'h2b15:	ff_dbi <= 8'h00;
		14'h2b16:	ff_dbi <= 8'h00;
		14'h2b17:	ff_dbi <= 8'h00;
		14'h2b18:	ff_dbi <= 8'h00;
		14'h2b19:	ff_dbi <= 8'h00;
		14'h2b1a:	ff_dbi <= 8'h00;
		14'h2b1b:	ff_dbi <= 8'h00;
		14'h2b1c:	ff_dbi <= 8'h00;
		14'h2b1d:	ff_dbi <= 8'h00;
		14'h2b1e:	ff_dbi <= 8'h00;
		14'h2b1f:	ff_dbi <= 8'h00;
		14'h2b20:	ff_dbi <= 8'h00;
		14'h2b21:	ff_dbi <= 8'h00;
		14'h2b22:	ff_dbi <= 8'h00;
		14'h2b23:	ff_dbi <= 8'h00;
		14'h2b24:	ff_dbi <= 8'h00;
		14'h2b25:	ff_dbi <= 8'h00;
		14'h2b26:	ff_dbi <= 8'h00;
		14'h2b27:	ff_dbi <= 8'h00;
		14'h2b28:	ff_dbi <= 8'h00;
		14'h2b29:	ff_dbi <= 8'h00;
		14'h2b2a:	ff_dbi <= 8'h00;
		14'h2b2b:	ff_dbi <= 8'h00;
		14'h2b2c:	ff_dbi <= 8'h00;
		14'h2b2d:	ff_dbi <= 8'h00;
		14'h2b2e:	ff_dbi <= 8'h00;
		14'h2b2f:	ff_dbi <= 8'h00;
		14'h2b30:	ff_dbi <= 8'h00;
		14'h2b31:	ff_dbi <= 8'h00;
		14'h2b32:	ff_dbi <= 8'h00;
		14'h2b33:	ff_dbi <= 8'h00;
		14'h2b34:	ff_dbi <= 8'h00;
		14'h2b35:	ff_dbi <= 8'h00;
		14'h2b36:	ff_dbi <= 8'h00;
		14'h2b37:	ff_dbi <= 8'h00;
		14'h2b38:	ff_dbi <= 8'h00;
		14'h2b39:	ff_dbi <= 8'h00;
		14'h2b3a:	ff_dbi <= 8'h00;
		14'h2b3b:	ff_dbi <= 8'h00;
		14'h2b3c:	ff_dbi <= 8'h00;
		14'h2b3d:	ff_dbi <= 8'h00;
		14'h2b3e:	ff_dbi <= 8'h00;
		14'h2b3f:	ff_dbi <= 8'h00;
		14'h2b40:	ff_dbi <= 8'h00;
		14'h2b41:	ff_dbi <= 8'h00;
		14'h2b42:	ff_dbi <= 8'h00;
		14'h2b43:	ff_dbi <= 8'h00;
		14'h2b44:	ff_dbi <= 8'h00;
		14'h2b45:	ff_dbi <= 8'h00;
		14'h2b46:	ff_dbi <= 8'h00;
		14'h2b47:	ff_dbi <= 8'h00;
		14'h2b48:	ff_dbi <= 8'h00;
		14'h2b49:	ff_dbi <= 8'h00;
		14'h2b4a:	ff_dbi <= 8'h00;
		14'h2b4b:	ff_dbi <= 8'h00;
		14'h2b4c:	ff_dbi <= 8'h00;
		14'h2b4d:	ff_dbi <= 8'h00;
		14'h2b4e:	ff_dbi <= 8'h00;
		14'h2b4f:	ff_dbi <= 8'h00;
		14'h2b50:	ff_dbi <= 8'h00;
		14'h2b51:	ff_dbi <= 8'h00;
		14'h2b52:	ff_dbi <= 8'h00;
		14'h2b53:	ff_dbi <= 8'h00;
		14'h2b54:	ff_dbi <= 8'h00;
		14'h2b55:	ff_dbi <= 8'h00;
		14'h2b56:	ff_dbi <= 8'h00;
		14'h2b57:	ff_dbi <= 8'h00;
		14'h2b58:	ff_dbi <= 8'h00;
		14'h2b59:	ff_dbi <= 8'h00;
		14'h2b5a:	ff_dbi <= 8'h00;
		14'h2b5b:	ff_dbi <= 8'h00;
		14'h2b5c:	ff_dbi <= 8'h00;
		14'h2b5d:	ff_dbi <= 8'h00;
		14'h2b5e:	ff_dbi <= 8'h00;
		14'h2b5f:	ff_dbi <= 8'h00;
		14'h2b60:	ff_dbi <= 8'h00;
		14'h2b61:	ff_dbi <= 8'h00;
		14'h2b62:	ff_dbi <= 8'h00;
		14'h2b63:	ff_dbi <= 8'h00;
		14'h2b64:	ff_dbi <= 8'h00;
		14'h2b65:	ff_dbi <= 8'h00;
		14'h2b66:	ff_dbi <= 8'h00;
		14'h2b67:	ff_dbi <= 8'h00;
		14'h2b68:	ff_dbi <= 8'h00;
		14'h2b69:	ff_dbi <= 8'h00;
		14'h2b6a:	ff_dbi <= 8'h00;
		14'h2b6b:	ff_dbi <= 8'h00;
		14'h2b6c:	ff_dbi <= 8'h00;
		14'h2b6d:	ff_dbi <= 8'h00;
		14'h2b6e:	ff_dbi <= 8'h00;
		14'h2b6f:	ff_dbi <= 8'h00;
		14'h2b70:	ff_dbi <= 8'h00;
		14'h2b71:	ff_dbi <= 8'h00;
		14'h2b72:	ff_dbi <= 8'h00;
		14'h2b73:	ff_dbi <= 8'h00;
		14'h2b74:	ff_dbi <= 8'h00;
		14'h2b75:	ff_dbi <= 8'h00;
		14'h2b76:	ff_dbi <= 8'h00;
		14'h2b77:	ff_dbi <= 8'h00;
		14'h2b78:	ff_dbi <= 8'h00;
		14'h2b79:	ff_dbi <= 8'h00;
		14'h2b7a:	ff_dbi <= 8'h00;
		14'h2b7b:	ff_dbi <= 8'h00;
		14'h2b7c:	ff_dbi <= 8'h00;
		14'h2b7d:	ff_dbi <= 8'h00;
		14'h2b7e:	ff_dbi <= 8'h00;
		14'h2b7f:	ff_dbi <= 8'h00;
		14'h2b80:	ff_dbi <= 8'h00;
		14'h2b81:	ff_dbi <= 8'h00;
		14'h2b82:	ff_dbi <= 8'h00;
		14'h2b83:	ff_dbi <= 8'h00;
		14'h2b84:	ff_dbi <= 8'h00;
		14'h2b85:	ff_dbi <= 8'h00;
		14'h2b86:	ff_dbi <= 8'h00;
		14'h2b87:	ff_dbi <= 8'h00;
		14'h2b88:	ff_dbi <= 8'h00;
		14'h2b89:	ff_dbi <= 8'h00;
		14'h2b8a:	ff_dbi <= 8'h00;
		14'h2b8b:	ff_dbi <= 8'h00;
		14'h2b8c:	ff_dbi <= 8'h00;
		14'h2b8d:	ff_dbi <= 8'h00;
		14'h2b8e:	ff_dbi <= 8'h00;
		14'h2b8f:	ff_dbi <= 8'h00;
		14'h2b90:	ff_dbi <= 8'h00;
		14'h2b91:	ff_dbi <= 8'h00;
		14'h2b92:	ff_dbi <= 8'h00;
		14'h2b93:	ff_dbi <= 8'h00;
		14'h2b94:	ff_dbi <= 8'h00;
		14'h2b95:	ff_dbi <= 8'h00;
		14'h2b96:	ff_dbi <= 8'h00;
		14'h2b97:	ff_dbi <= 8'h00;
		14'h2b98:	ff_dbi <= 8'h00;
		14'h2b99:	ff_dbi <= 8'h00;
		14'h2b9a:	ff_dbi <= 8'h00;
		14'h2b9b:	ff_dbi <= 8'h00;
		14'h2b9c:	ff_dbi <= 8'h00;
		14'h2b9d:	ff_dbi <= 8'h00;
		14'h2b9e:	ff_dbi <= 8'h00;
		14'h2b9f:	ff_dbi <= 8'h00;
		14'h2ba0:	ff_dbi <= 8'h00;
		14'h2ba1:	ff_dbi <= 8'h00;
		14'h2ba2:	ff_dbi <= 8'h00;
		14'h2ba3:	ff_dbi <= 8'h00;
		14'h2ba4:	ff_dbi <= 8'h00;
		14'h2ba5:	ff_dbi <= 8'h00;
		14'h2ba6:	ff_dbi <= 8'h00;
		14'h2ba7:	ff_dbi <= 8'h00;
		14'h2ba8:	ff_dbi <= 8'h00;
		14'h2ba9:	ff_dbi <= 8'h00;
		14'h2baa:	ff_dbi <= 8'h00;
		14'h2bab:	ff_dbi <= 8'h00;
		14'h2bac:	ff_dbi <= 8'h00;
		14'h2bad:	ff_dbi <= 8'h00;
		14'h2bae:	ff_dbi <= 8'h00;
		14'h2baf:	ff_dbi <= 8'h00;
		14'h2bb0:	ff_dbi <= 8'h00;
		14'h2bb1:	ff_dbi <= 8'h00;
		14'h2bb2:	ff_dbi <= 8'h00;
		14'h2bb3:	ff_dbi <= 8'h00;
		14'h2bb4:	ff_dbi <= 8'h00;
		14'h2bb5:	ff_dbi <= 8'h00;
		14'h2bb6:	ff_dbi <= 8'h00;
		14'h2bb7:	ff_dbi <= 8'h00;
		14'h2bb8:	ff_dbi <= 8'h00;
		14'h2bb9:	ff_dbi <= 8'h00;
		14'h2bba:	ff_dbi <= 8'h00;
		14'h2bbb:	ff_dbi <= 8'h00;
		14'h2bbc:	ff_dbi <= 8'h00;
		14'h2bbd:	ff_dbi <= 8'h00;
		14'h2bbe:	ff_dbi <= 8'h00;
		14'h2bbf:	ff_dbi <= 8'h00;
		14'h2bc0:	ff_dbi <= 8'h00;
		14'h2bc1:	ff_dbi <= 8'h00;
		14'h2bc2:	ff_dbi <= 8'h00;
		14'h2bc3:	ff_dbi <= 8'h00;
		14'h2bc4:	ff_dbi <= 8'h00;
		14'h2bc5:	ff_dbi <= 8'h00;
		14'h2bc6:	ff_dbi <= 8'h00;
		14'h2bc7:	ff_dbi <= 8'h00;
		14'h2bc8:	ff_dbi <= 8'h00;
		14'h2bc9:	ff_dbi <= 8'h00;
		14'h2bca:	ff_dbi <= 8'h00;
		14'h2bcb:	ff_dbi <= 8'h00;
		14'h2bcc:	ff_dbi <= 8'h00;
		14'h2bcd:	ff_dbi <= 8'h00;
		14'h2bce:	ff_dbi <= 8'h00;
		14'h2bcf:	ff_dbi <= 8'h00;
		14'h2bd0:	ff_dbi <= 8'h00;
		14'h2bd1:	ff_dbi <= 8'h00;
		14'h2bd2:	ff_dbi <= 8'h00;
		14'h2bd3:	ff_dbi <= 8'h00;
		14'h2bd4:	ff_dbi <= 8'h00;
		14'h2bd5:	ff_dbi <= 8'h00;
		14'h2bd6:	ff_dbi <= 8'h00;
		14'h2bd7:	ff_dbi <= 8'h00;
		14'h2bd8:	ff_dbi <= 8'h00;
		14'h2bd9:	ff_dbi <= 8'h00;
		14'h2bda:	ff_dbi <= 8'h00;
		14'h2bdb:	ff_dbi <= 8'h00;
		14'h2bdc:	ff_dbi <= 8'h00;
		14'h2bdd:	ff_dbi <= 8'h00;
		14'h2bde:	ff_dbi <= 8'h00;
		14'h2bdf:	ff_dbi <= 8'h00;
		14'h2be0:	ff_dbi <= 8'h00;
		14'h2be1:	ff_dbi <= 8'h00;
		14'h2be2:	ff_dbi <= 8'h00;
		14'h2be3:	ff_dbi <= 8'h00;
		14'h2be4:	ff_dbi <= 8'h00;
		14'h2be5:	ff_dbi <= 8'h00;
		14'h2be6:	ff_dbi <= 8'h00;
		14'h2be7:	ff_dbi <= 8'h00;
		14'h2be8:	ff_dbi <= 8'h00;
		14'h2be9:	ff_dbi <= 8'h00;
		14'h2bea:	ff_dbi <= 8'h00;
		14'h2beb:	ff_dbi <= 8'h00;
		14'h2bec:	ff_dbi <= 8'h00;
		14'h2bed:	ff_dbi <= 8'h00;
		14'h2bee:	ff_dbi <= 8'h00;
		14'h2bef:	ff_dbi <= 8'h00;
		14'h2bf0:	ff_dbi <= 8'h00;
		14'h2bf1:	ff_dbi <= 8'h00;
		14'h2bf2:	ff_dbi <= 8'h00;
		14'h2bf3:	ff_dbi <= 8'h00;
		14'h2bf4:	ff_dbi <= 8'h00;
		14'h2bf5:	ff_dbi <= 8'h00;
		14'h2bf6:	ff_dbi <= 8'h00;
		14'h2bf7:	ff_dbi <= 8'h00;
		14'h2bf8:	ff_dbi <= 8'h00;
		14'h2bf9:	ff_dbi <= 8'h00;
		14'h2bfa:	ff_dbi <= 8'h00;
		14'h2bfb:	ff_dbi <= 8'h00;
		14'h2bfc:	ff_dbi <= 8'h00;
		14'h2bfd:	ff_dbi <= 8'h00;
		14'h2bfe:	ff_dbi <= 8'h00;
		14'h2bff:	ff_dbi <= 8'h00;
		14'h2c00:	ff_dbi <= 8'h00;
		14'h2c01:	ff_dbi <= 8'h00;
		14'h2c02:	ff_dbi <= 8'h00;
		14'h2c03:	ff_dbi <= 8'h00;
		14'h2c04:	ff_dbi <= 8'h00;
		14'h2c05:	ff_dbi <= 8'h00;
		14'h2c06:	ff_dbi <= 8'h00;
		14'h2c07:	ff_dbi <= 8'h00;
		14'h2c08:	ff_dbi <= 8'h00;
		14'h2c09:	ff_dbi <= 8'h00;
		14'h2c0a:	ff_dbi <= 8'h00;
		14'h2c0b:	ff_dbi <= 8'h00;
		14'h2c0c:	ff_dbi <= 8'h00;
		14'h2c0d:	ff_dbi <= 8'h00;
		14'h2c0e:	ff_dbi <= 8'h00;
		14'h2c0f:	ff_dbi <= 8'h00;
		14'h2c10:	ff_dbi <= 8'h00;
		14'h2c11:	ff_dbi <= 8'h00;
		14'h2c12:	ff_dbi <= 8'h00;
		14'h2c13:	ff_dbi <= 8'h00;
		14'h2c14:	ff_dbi <= 8'h00;
		14'h2c15:	ff_dbi <= 8'h00;
		14'h2c16:	ff_dbi <= 8'h00;
		14'h2c17:	ff_dbi <= 8'h00;
		14'h2c18:	ff_dbi <= 8'h00;
		14'h2c19:	ff_dbi <= 8'h00;
		14'h2c1a:	ff_dbi <= 8'h00;
		14'h2c1b:	ff_dbi <= 8'h00;
		14'h2c1c:	ff_dbi <= 8'h00;
		14'h2c1d:	ff_dbi <= 8'h00;
		14'h2c1e:	ff_dbi <= 8'h00;
		14'h2c1f:	ff_dbi <= 8'h00;
		14'h2c20:	ff_dbi <= 8'h00;
		14'h2c21:	ff_dbi <= 8'h00;
		14'h2c22:	ff_dbi <= 8'h00;
		14'h2c23:	ff_dbi <= 8'h00;
		14'h2c24:	ff_dbi <= 8'h00;
		14'h2c25:	ff_dbi <= 8'h00;
		14'h2c26:	ff_dbi <= 8'h00;
		14'h2c27:	ff_dbi <= 8'h00;
		14'h2c28:	ff_dbi <= 8'h00;
		14'h2c29:	ff_dbi <= 8'h00;
		14'h2c2a:	ff_dbi <= 8'h00;
		14'h2c2b:	ff_dbi <= 8'h00;
		14'h2c2c:	ff_dbi <= 8'h00;
		14'h2c2d:	ff_dbi <= 8'h00;
		14'h2c2e:	ff_dbi <= 8'h00;
		14'h2c2f:	ff_dbi <= 8'h00;
		14'h2c30:	ff_dbi <= 8'h00;
		14'h2c31:	ff_dbi <= 8'h00;
		14'h2c32:	ff_dbi <= 8'h00;
		14'h2c33:	ff_dbi <= 8'h00;
		14'h2c34:	ff_dbi <= 8'h00;
		14'h2c35:	ff_dbi <= 8'h00;
		14'h2c36:	ff_dbi <= 8'h00;
		14'h2c37:	ff_dbi <= 8'h00;
		14'h2c38:	ff_dbi <= 8'h00;
		14'h2c39:	ff_dbi <= 8'h00;
		14'h2c3a:	ff_dbi <= 8'h00;
		14'h2c3b:	ff_dbi <= 8'h00;
		14'h2c3c:	ff_dbi <= 8'h00;
		14'h2c3d:	ff_dbi <= 8'h00;
		14'h2c3e:	ff_dbi <= 8'h00;
		14'h2c3f:	ff_dbi <= 8'h00;
		14'h2c40:	ff_dbi <= 8'h00;
		14'h2c41:	ff_dbi <= 8'h00;
		14'h2c42:	ff_dbi <= 8'h00;
		14'h2c43:	ff_dbi <= 8'h00;
		14'h2c44:	ff_dbi <= 8'h00;
		14'h2c45:	ff_dbi <= 8'h00;
		14'h2c46:	ff_dbi <= 8'h00;
		14'h2c47:	ff_dbi <= 8'h00;
		14'h2c48:	ff_dbi <= 8'h00;
		14'h2c49:	ff_dbi <= 8'h00;
		14'h2c4a:	ff_dbi <= 8'h00;
		14'h2c4b:	ff_dbi <= 8'h00;
		14'h2c4c:	ff_dbi <= 8'h00;
		14'h2c4d:	ff_dbi <= 8'h00;
		14'h2c4e:	ff_dbi <= 8'h00;
		14'h2c4f:	ff_dbi <= 8'h00;
		14'h2c50:	ff_dbi <= 8'h00;
		14'h2c51:	ff_dbi <= 8'h00;
		14'h2c52:	ff_dbi <= 8'h00;
		14'h2c53:	ff_dbi <= 8'h00;
		14'h2c54:	ff_dbi <= 8'h00;
		14'h2c55:	ff_dbi <= 8'h00;
		14'h2c56:	ff_dbi <= 8'h00;
		14'h2c57:	ff_dbi <= 8'h00;
		14'h2c58:	ff_dbi <= 8'h00;
		14'h2c59:	ff_dbi <= 8'h00;
		14'h2c5a:	ff_dbi <= 8'h00;
		14'h2c5b:	ff_dbi <= 8'h00;
		14'h2c5c:	ff_dbi <= 8'h00;
		14'h2c5d:	ff_dbi <= 8'h00;
		14'h2c5e:	ff_dbi <= 8'h00;
		14'h2c5f:	ff_dbi <= 8'h00;
		14'h2c60:	ff_dbi <= 8'h00;
		14'h2c61:	ff_dbi <= 8'h00;
		14'h2c62:	ff_dbi <= 8'h00;
		14'h2c63:	ff_dbi <= 8'h00;
		14'h2c64:	ff_dbi <= 8'h00;
		14'h2c65:	ff_dbi <= 8'h00;
		14'h2c66:	ff_dbi <= 8'h00;
		14'h2c67:	ff_dbi <= 8'h00;
		14'h2c68:	ff_dbi <= 8'h00;
		14'h2c69:	ff_dbi <= 8'h00;
		14'h2c6a:	ff_dbi <= 8'h00;
		14'h2c6b:	ff_dbi <= 8'h00;
		14'h2c6c:	ff_dbi <= 8'h00;
		14'h2c6d:	ff_dbi <= 8'h00;
		14'h2c6e:	ff_dbi <= 8'h00;
		14'h2c6f:	ff_dbi <= 8'h00;
		14'h2c70:	ff_dbi <= 8'h00;
		14'h2c71:	ff_dbi <= 8'h00;
		14'h2c72:	ff_dbi <= 8'h00;
		14'h2c73:	ff_dbi <= 8'h00;
		14'h2c74:	ff_dbi <= 8'h00;
		14'h2c75:	ff_dbi <= 8'h00;
		14'h2c76:	ff_dbi <= 8'h00;
		14'h2c77:	ff_dbi <= 8'h00;
		14'h2c78:	ff_dbi <= 8'h00;
		14'h2c79:	ff_dbi <= 8'h00;
		14'h2c7a:	ff_dbi <= 8'h00;
		14'h2c7b:	ff_dbi <= 8'h00;
		14'h2c7c:	ff_dbi <= 8'h00;
		14'h2c7d:	ff_dbi <= 8'h00;
		14'h2c7e:	ff_dbi <= 8'h00;
		14'h2c7f:	ff_dbi <= 8'h00;
		14'h2c80:	ff_dbi <= 8'h00;
		14'h2c81:	ff_dbi <= 8'h00;
		14'h2c82:	ff_dbi <= 8'h00;
		14'h2c83:	ff_dbi <= 8'h00;
		14'h2c84:	ff_dbi <= 8'h00;
		14'h2c85:	ff_dbi <= 8'h00;
		14'h2c86:	ff_dbi <= 8'h00;
		14'h2c87:	ff_dbi <= 8'h00;
		14'h2c88:	ff_dbi <= 8'h00;
		14'h2c89:	ff_dbi <= 8'h00;
		14'h2c8a:	ff_dbi <= 8'h00;
		14'h2c8b:	ff_dbi <= 8'h00;
		14'h2c8c:	ff_dbi <= 8'h00;
		14'h2c8d:	ff_dbi <= 8'h00;
		14'h2c8e:	ff_dbi <= 8'h00;
		14'h2c8f:	ff_dbi <= 8'h00;
		14'h2c90:	ff_dbi <= 8'h00;
		14'h2c91:	ff_dbi <= 8'h00;
		14'h2c92:	ff_dbi <= 8'h00;
		14'h2c93:	ff_dbi <= 8'h00;
		14'h2c94:	ff_dbi <= 8'h00;
		14'h2c95:	ff_dbi <= 8'h00;
		14'h2c96:	ff_dbi <= 8'h00;
		14'h2c97:	ff_dbi <= 8'h00;
		14'h2c98:	ff_dbi <= 8'h00;
		14'h2c99:	ff_dbi <= 8'h00;
		14'h2c9a:	ff_dbi <= 8'h00;
		14'h2c9b:	ff_dbi <= 8'h00;
		14'h2c9c:	ff_dbi <= 8'h00;
		14'h2c9d:	ff_dbi <= 8'h00;
		14'h2c9e:	ff_dbi <= 8'h00;
		14'h2c9f:	ff_dbi <= 8'h00;
		14'h2ca0:	ff_dbi <= 8'h00;
		14'h2ca1:	ff_dbi <= 8'h00;
		14'h2ca2:	ff_dbi <= 8'h00;
		14'h2ca3:	ff_dbi <= 8'h00;
		14'h2ca4:	ff_dbi <= 8'h00;
		14'h2ca5:	ff_dbi <= 8'h00;
		14'h2ca6:	ff_dbi <= 8'h00;
		14'h2ca7:	ff_dbi <= 8'h00;
		14'h2ca8:	ff_dbi <= 8'h00;
		14'h2ca9:	ff_dbi <= 8'h00;
		14'h2caa:	ff_dbi <= 8'h00;
		14'h2cab:	ff_dbi <= 8'h00;
		14'h2cac:	ff_dbi <= 8'h00;
		14'h2cad:	ff_dbi <= 8'h00;
		14'h2cae:	ff_dbi <= 8'h00;
		14'h2caf:	ff_dbi <= 8'h00;
		14'h2cb0:	ff_dbi <= 8'h00;
		14'h2cb1:	ff_dbi <= 8'h00;
		14'h2cb2:	ff_dbi <= 8'h00;
		14'h2cb3:	ff_dbi <= 8'h00;
		14'h2cb4:	ff_dbi <= 8'h00;
		14'h2cb5:	ff_dbi <= 8'h00;
		14'h2cb6:	ff_dbi <= 8'h00;
		14'h2cb7:	ff_dbi <= 8'h00;
		14'h2cb8:	ff_dbi <= 8'h00;
		14'h2cb9:	ff_dbi <= 8'h00;
		14'h2cba:	ff_dbi <= 8'h00;
		14'h2cbb:	ff_dbi <= 8'h00;
		14'h2cbc:	ff_dbi <= 8'h00;
		14'h2cbd:	ff_dbi <= 8'h00;
		14'h2cbe:	ff_dbi <= 8'h00;
		14'h2cbf:	ff_dbi <= 8'h00;
		14'h2cc0:	ff_dbi <= 8'h00;
		14'h2cc1:	ff_dbi <= 8'h00;
		14'h2cc2:	ff_dbi <= 8'h00;
		14'h2cc3:	ff_dbi <= 8'h00;
		14'h2cc4:	ff_dbi <= 8'h00;
		14'h2cc5:	ff_dbi <= 8'h00;
		14'h2cc6:	ff_dbi <= 8'h00;
		14'h2cc7:	ff_dbi <= 8'h00;
		14'h2cc8:	ff_dbi <= 8'h00;
		14'h2cc9:	ff_dbi <= 8'h00;
		14'h2cca:	ff_dbi <= 8'h00;
		14'h2ccb:	ff_dbi <= 8'h00;
		14'h2ccc:	ff_dbi <= 8'h00;
		14'h2ccd:	ff_dbi <= 8'h00;
		14'h2cce:	ff_dbi <= 8'h00;
		14'h2ccf:	ff_dbi <= 8'h00;
		14'h2cd0:	ff_dbi <= 8'h00;
		14'h2cd1:	ff_dbi <= 8'h00;
		14'h2cd2:	ff_dbi <= 8'h00;
		14'h2cd3:	ff_dbi <= 8'h00;
		14'h2cd4:	ff_dbi <= 8'h00;
		14'h2cd5:	ff_dbi <= 8'h00;
		14'h2cd6:	ff_dbi <= 8'h00;
		14'h2cd7:	ff_dbi <= 8'h00;
		14'h2cd8:	ff_dbi <= 8'h00;
		14'h2cd9:	ff_dbi <= 8'h00;
		14'h2cda:	ff_dbi <= 8'h00;
		14'h2cdb:	ff_dbi <= 8'h00;
		14'h2cdc:	ff_dbi <= 8'h00;
		14'h2cdd:	ff_dbi <= 8'h00;
		14'h2cde:	ff_dbi <= 8'h00;
		14'h2cdf:	ff_dbi <= 8'h00;
		14'h2ce0:	ff_dbi <= 8'h00;
		14'h2ce1:	ff_dbi <= 8'h00;
		14'h2ce2:	ff_dbi <= 8'h00;
		14'h2ce3:	ff_dbi <= 8'h00;
		14'h2ce4:	ff_dbi <= 8'h00;
		14'h2ce5:	ff_dbi <= 8'h00;
		14'h2ce6:	ff_dbi <= 8'h00;
		14'h2ce7:	ff_dbi <= 8'h00;
		14'h2ce8:	ff_dbi <= 8'h00;
		14'h2ce9:	ff_dbi <= 8'h00;
		14'h2cea:	ff_dbi <= 8'h00;
		14'h2ceb:	ff_dbi <= 8'h00;
		14'h2cec:	ff_dbi <= 8'h00;
		14'h2ced:	ff_dbi <= 8'h00;
		14'h2cee:	ff_dbi <= 8'h00;
		14'h2cef:	ff_dbi <= 8'h00;
		14'h2cf0:	ff_dbi <= 8'h00;
		14'h2cf1:	ff_dbi <= 8'h00;
		14'h2cf2:	ff_dbi <= 8'h00;
		14'h2cf3:	ff_dbi <= 8'h00;
		14'h2cf4:	ff_dbi <= 8'h00;
		14'h2cf5:	ff_dbi <= 8'h00;
		14'h2cf6:	ff_dbi <= 8'h00;
		14'h2cf7:	ff_dbi <= 8'h00;
		14'h2cf8:	ff_dbi <= 8'h00;
		14'h2cf9:	ff_dbi <= 8'h00;
		14'h2cfa:	ff_dbi <= 8'h00;
		14'h2cfb:	ff_dbi <= 8'h00;
		14'h2cfc:	ff_dbi <= 8'h00;
		14'h2cfd:	ff_dbi <= 8'h00;
		14'h2cfe:	ff_dbi <= 8'h00;
		14'h2cff:	ff_dbi <= 8'h00;
		14'h2d00:	ff_dbi <= 8'h00;
		14'h2d01:	ff_dbi <= 8'h00;
		14'h2d02:	ff_dbi <= 8'h00;
		14'h2d03:	ff_dbi <= 8'h00;
		14'h2d04:	ff_dbi <= 8'h00;
		14'h2d05:	ff_dbi <= 8'h00;
		14'h2d06:	ff_dbi <= 8'h00;
		14'h2d07:	ff_dbi <= 8'h00;
		14'h2d08:	ff_dbi <= 8'h00;
		14'h2d09:	ff_dbi <= 8'h00;
		14'h2d0a:	ff_dbi <= 8'h00;
		14'h2d0b:	ff_dbi <= 8'h00;
		14'h2d0c:	ff_dbi <= 8'h00;
		14'h2d0d:	ff_dbi <= 8'h00;
		14'h2d0e:	ff_dbi <= 8'h00;
		14'h2d0f:	ff_dbi <= 8'h00;
		14'h2d10:	ff_dbi <= 8'h00;
		14'h2d11:	ff_dbi <= 8'h00;
		14'h2d12:	ff_dbi <= 8'h00;
		14'h2d13:	ff_dbi <= 8'h00;
		14'h2d14:	ff_dbi <= 8'h00;
		14'h2d15:	ff_dbi <= 8'h00;
		14'h2d16:	ff_dbi <= 8'h00;
		14'h2d17:	ff_dbi <= 8'h00;
		14'h2d18:	ff_dbi <= 8'h00;
		14'h2d19:	ff_dbi <= 8'h00;
		14'h2d1a:	ff_dbi <= 8'h00;
		14'h2d1b:	ff_dbi <= 8'h00;
		14'h2d1c:	ff_dbi <= 8'h00;
		14'h2d1d:	ff_dbi <= 8'h00;
		14'h2d1e:	ff_dbi <= 8'h00;
		14'h2d1f:	ff_dbi <= 8'h00;
		14'h2d20:	ff_dbi <= 8'h00;
		14'h2d21:	ff_dbi <= 8'h00;
		14'h2d22:	ff_dbi <= 8'h00;
		14'h2d23:	ff_dbi <= 8'h00;
		14'h2d24:	ff_dbi <= 8'h00;
		14'h2d25:	ff_dbi <= 8'h00;
		14'h2d26:	ff_dbi <= 8'h00;
		14'h2d27:	ff_dbi <= 8'h00;
		14'h2d28:	ff_dbi <= 8'h00;
		14'h2d29:	ff_dbi <= 8'h00;
		14'h2d2a:	ff_dbi <= 8'h00;
		14'h2d2b:	ff_dbi <= 8'h00;
		14'h2d2c:	ff_dbi <= 8'h00;
		14'h2d2d:	ff_dbi <= 8'h00;
		14'h2d2e:	ff_dbi <= 8'h00;
		14'h2d2f:	ff_dbi <= 8'h00;
		14'h2d30:	ff_dbi <= 8'h00;
		14'h2d31:	ff_dbi <= 8'h00;
		14'h2d32:	ff_dbi <= 8'h00;
		14'h2d33:	ff_dbi <= 8'h00;
		14'h2d34:	ff_dbi <= 8'h00;
		14'h2d35:	ff_dbi <= 8'h00;
		14'h2d36:	ff_dbi <= 8'h00;
		14'h2d37:	ff_dbi <= 8'h00;
		14'h2d38:	ff_dbi <= 8'h00;
		14'h2d39:	ff_dbi <= 8'h00;
		14'h2d3a:	ff_dbi <= 8'h00;
		14'h2d3b:	ff_dbi <= 8'h00;
		14'h2d3c:	ff_dbi <= 8'h00;
		14'h2d3d:	ff_dbi <= 8'h00;
		14'h2d3e:	ff_dbi <= 8'h00;
		14'h2d3f:	ff_dbi <= 8'h00;
		14'h2d40:	ff_dbi <= 8'h00;
		14'h2d41:	ff_dbi <= 8'h00;
		14'h2d42:	ff_dbi <= 8'h00;
		14'h2d43:	ff_dbi <= 8'h00;
		14'h2d44:	ff_dbi <= 8'h00;
		14'h2d45:	ff_dbi <= 8'h00;
		14'h2d46:	ff_dbi <= 8'h00;
		14'h2d47:	ff_dbi <= 8'h00;
		14'h2d48:	ff_dbi <= 8'h00;
		14'h2d49:	ff_dbi <= 8'h00;
		14'h2d4a:	ff_dbi <= 8'h00;
		14'h2d4b:	ff_dbi <= 8'h00;
		14'h2d4c:	ff_dbi <= 8'h00;
		14'h2d4d:	ff_dbi <= 8'h00;
		14'h2d4e:	ff_dbi <= 8'h00;
		14'h2d4f:	ff_dbi <= 8'h00;
		14'h2d50:	ff_dbi <= 8'h00;
		14'h2d51:	ff_dbi <= 8'h00;
		14'h2d52:	ff_dbi <= 8'h00;
		14'h2d53:	ff_dbi <= 8'h00;
		14'h2d54:	ff_dbi <= 8'h00;
		14'h2d55:	ff_dbi <= 8'h00;
		14'h2d56:	ff_dbi <= 8'h00;
		14'h2d57:	ff_dbi <= 8'h00;
		14'h2d58:	ff_dbi <= 8'h00;
		14'h2d59:	ff_dbi <= 8'h00;
		14'h2d5a:	ff_dbi <= 8'h00;
		14'h2d5b:	ff_dbi <= 8'h00;
		14'h2d5c:	ff_dbi <= 8'h00;
		14'h2d5d:	ff_dbi <= 8'h00;
		14'h2d5e:	ff_dbi <= 8'h00;
		14'h2d5f:	ff_dbi <= 8'h00;
		14'h2d60:	ff_dbi <= 8'h00;
		14'h2d61:	ff_dbi <= 8'h00;
		14'h2d62:	ff_dbi <= 8'h00;
		14'h2d63:	ff_dbi <= 8'h00;
		14'h2d64:	ff_dbi <= 8'h00;
		14'h2d65:	ff_dbi <= 8'h00;
		14'h2d66:	ff_dbi <= 8'h00;
		14'h2d67:	ff_dbi <= 8'h00;
		14'h2d68:	ff_dbi <= 8'h00;
		14'h2d69:	ff_dbi <= 8'h00;
		14'h2d6a:	ff_dbi <= 8'h00;
		14'h2d6b:	ff_dbi <= 8'h00;
		14'h2d6c:	ff_dbi <= 8'h00;
		14'h2d6d:	ff_dbi <= 8'h00;
		14'h2d6e:	ff_dbi <= 8'h00;
		14'h2d6f:	ff_dbi <= 8'h00;
		14'h2d70:	ff_dbi <= 8'h00;
		14'h2d71:	ff_dbi <= 8'h00;
		14'h2d72:	ff_dbi <= 8'h00;
		14'h2d73:	ff_dbi <= 8'h00;
		14'h2d74:	ff_dbi <= 8'h00;
		14'h2d75:	ff_dbi <= 8'h00;
		14'h2d76:	ff_dbi <= 8'h00;
		14'h2d77:	ff_dbi <= 8'h00;
		14'h2d78:	ff_dbi <= 8'h00;
		14'h2d79:	ff_dbi <= 8'h00;
		14'h2d7a:	ff_dbi <= 8'h00;
		14'h2d7b:	ff_dbi <= 8'h00;
		14'h2d7c:	ff_dbi <= 8'h00;
		14'h2d7d:	ff_dbi <= 8'h00;
		14'h2d7e:	ff_dbi <= 8'h00;
		14'h2d7f:	ff_dbi <= 8'h00;
		14'h2d80:	ff_dbi <= 8'h00;
		14'h2d81:	ff_dbi <= 8'h00;
		14'h2d82:	ff_dbi <= 8'h00;
		14'h2d83:	ff_dbi <= 8'h00;
		14'h2d84:	ff_dbi <= 8'h00;
		14'h2d85:	ff_dbi <= 8'h00;
		14'h2d86:	ff_dbi <= 8'h00;
		14'h2d87:	ff_dbi <= 8'h00;
		14'h2d88:	ff_dbi <= 8'h00;
		14'h2d89:	ff_dbi <= 8'h00;
		14'h2d8a:	ff_dbi <= 8'h00;
		14'h2d8b:	ff_dbi <= 8'h00;
		14'h2d8c:	ff_dbi <= 8'h00;
		14'h2d8d:	ff_dbi <= 8'h00;
		14'h2d8e:	ff_dbi <= 8'h00;
		14'h2d8f:	ff_dbi <= 8'h00;
		14'h2d90:	ff_dbi <= 8'h00;
		14'h2d91:	ff_dbi <= 8'h00;
		14'h2d92:	ff_dbi <= 8'h00;
		14'h2d93:	ff_dbi <= 8'h00;
		14'h2d94:	ff_dbi <= 8'h00;
		14'h2d95:	ff_dbi <= 8'h00;
		14'h2d96:	ff_dbi <= 8'h00;
		14'h2d97:	ff_dbi <= 8'h00;
		14'h2d98:	ff_dbi <= 8'h00;
		14'h2d99:	ff_dbi <= 8'h00;
		14'h2d9a:	ff_dbi <= 8'h00;
		14'h2d9b:	ff_dbi <= 8'h00;
		14'h2d9c:	ff_dbi <= 8'h00;
		14'h2d9d:	ff_dbi <= 8'h00;
		14'h2d9e:	ff_dbi <= 8'h00;
		14'h2d9f:	ff_dbi <= 8'h00;
		14'h2da0:	ff_dbi <= 8'h00;
		14'h2da1:	ff_dbi <= 8'h00;
		14'h2da2:	ff_dbi <= 8'h00;
		14'h2da3:	ff_dbi <= 8'h00;
		14'h2da4:	ff_dbi <= 8'h00;
		14'h2da5:	ff_dbi <= 8'h00;
		14'h2da6:	ff_dbi <= 8'h00;
		14'h2da7:	ff_dbi <= 8'h00;
		14'h2da8:	ff_dbi <= 8'h00;
		14'h2da9:	ff_dbi <= 8'h00;
		14'h2daa:	ff_dbi <= 8'h00;
		14'h2dab:	ff_dbi <= 8'h00;
		14'h2dac:	ff_dbi <= 8'h00;
		14'h2dad:	ff_dbi <= 8'h00;
		14'h2dae:	ff_dbi <= 8'h00;
		14'h2daf:	ff_dbi <= 8'h00;
		14'h2db0:	ff_dbi <= 8'h00;
		14'h2db1:	ff_dbi <= 8'h00;
		14'h2db2:	ff_dbi <= 8'h00;
		14'h2db3:	ff_dbi <= 8'h00;
		14'h2db4:	ff_dbi <= 8'h00;
		14'h2db5:	ff_dbi <= 8'h00;
		14'h2db6:	ff_dbi <= 8'h00;
		14'h2db7:	ff_dbi <= 8'h00;
		14'h2db8:	ff_dbi <= 8'h00;
		14'h2db9:	ff_dbi <= 8'h00;
		14'h2dba:	ff_dbi <= 8'h00;
		14'h2dbb:	ff_dbi <= 8'h00;
		14'h2dbc:	ff_dbi <= 8'h00;
		14'h2dbd:	ff_dbi <= 8'h00;
		14'h2dbe:	ff_dbi <= 8'h00;
		14'h2dbf:	ff_dbi <= 8'h00;
		14'h2dc0:	ff_dbi <= 8'h00;
		14'h2dc1:	ff_dbi <= 8'h00;
		14'h2dc2:	ff_dbi <= 8'h00;
		14'h2dc3:	ff_dbi <= 8'h00;
		14'h2dc4:	ff_dbi <= 8'h00;
		14'h2dc5:	ff_dbi <= 8'h00;
		14'h2dc6:	ff_dbi <= 8'h00;
		14'h2dc7:	ff_dbi <= 8'h00;
		14'h2dc8:	ff_dbi <= 8'h00;
		14'h2dc9:	ff_dbi <= 8'h00;
		14'h2dca:	ff_dbi <= 8'h00;
		14'h2dcb:	ff_dbi <= 8'h00;
		14'h2dcc:	ff_dbi <= 8'h00;
		14'h2dcd:	ff_dbi <= 8'h00;
		14'h2dce:	ff_dbi <= 8'h00;
		14'h2dcf:	ff_dbi <= 8'h00;
		14'h2dd0:	ff_dbi <= 8'h00;
		14'h2dd1:	ff_dbi <= 8'h00;
		14'h2dd2:	ff_dbi <= 8'h00;
		14'h2dd3:	ff_dbi <= 8'h00;
		14'h2dd4:	ff_dbi <= 8'h00;
		14'h2dd5:	ff_dbi <= 8'h00;
		14'h2dd6:	ff_dbi <= 8'h00;
		14'h2dd7:	ff_dbi <= 8'h00;
		14'h2dd8:	ff_dbi <= 8'h00;
		14'h2dd9:	ff_dbi <= 8'h00;
		14'h2dda:	ff_dbi <= 8'h00;
		14'h2ddb:	ff_dbi <= 8'h00;
		14'h2ddc:	ff_dbi <= 8'h00;
		14'h2ddd:	ff_dbi <= 8'h00;
		14'h2dde:	ff_dbi <= 8'h00;
		14'h2ddf:	ff_dbi <= 8'h00;
		14'h2de0:	ff_dbi <= 8'h00;
		14'h2de1:	ff_dbi <= 8'h00;
		14'h2de2:	ff_dbi <= 8'h00;
		14'h2de3:	ff_dbi <= 8'h00;
		14'h2de4:	ff_dbi <= 8'h00;
		14'h2de5:	ff_dbi <= 8'h00;
		14'h2de6:	ff_dbi <= 8'h00;
		14'h2de7:	ff_dbi <= 8'h00;
		14'h2de8:	ff_dbi <= 8'h00;
		14'h2de9:	ff_dbi <= 8'h00;
		14'h2dea:	ff_dbi <= 8'h00;
		14'h2deb:	ff_dbi <= 8'h00;
		14'h2dec:	ff_dbi <= 8'h00;
		14'h2ded:	ff_dbi <= 8'h00;
		14'h2dee:	ff_dbi <= 8'h00;
		14'h2def:	ff_dbi <= 8'h00;
		14'h2df0:	ff_dbi <= 8'h00;
		14'h2df1:	ff_dbi <= 8'h00;
		14'h2df2:	ff_dbi <= 8'h00;
		14'h2df3:	ff_dbi <= 8'h00;
		14'h2df4:	ff_dbi <= 8'h00;
		14'h2df5:	ff_dbi <= 8'h00;
		14'h2df6:	ff_dbi <= 8'h00;
		14'h2df7:	ff_dbi <= 8'h00;
		14'h2df8:	ff_dbi <= 8'h00;
		14'h2df9:	ff_dbi <= 8'h00;
		14'h2dfa:	ff_dbi <= 8'h00;
		14'h2dfb:	ff_dbi <= 8'h00;
		14'h2dfc:	ff_dbi <= 8'h00;
		14'h2dfd:	ff_dbi <= 8'h00;
		14'h2dfe:	ff_dbi <= 8'h00;
		14'h2dff:	ff_dbi <= 8'h00;
		14'h2e00:	ff_dbi <= 8'h00;
		14'h2e01:	ff_dbi <= 8'h00;
		14'h2e02:	ff_dbi <= 8'h00;
		14'h2e03:	ff_dbi <= 8'h00;
		14'h2e04:	ff_dbi <= 8'h00;
		14'h2e05:	ff_dbi <= 8'h00;
		14'h2e06:	ff_dbi <= 8'h00;
		14'h2e07:	ff_dbi <= 8'h00;
		14'h2e08:	ff_dbi <= 8'h00;
		14'h2e09:	ff_dbi <= 8'h00;
		14'h2e0a:	ff_dbi <= 8'h00;
		14'h2e0b:	ff_dbi <= 8'h00;
		14'h2e0c:	ff_dbi <= 8'h00;
		14'h2e0d:	ff_dbi <= 8'h00;
		14'h2e0e:	ff_dbi <= 8'h00;
		14'h2e0f:	ff_dbi <= 8'h00;
		14'h2e10:	ff_dbi <= 8'h00;
		14'h2e11:	ff_dbi <= 8'h00;
		14'h2e12:	ff_dbi <= 8'h00;
		14'h2e13:	ff_dbi <= 8'h00;
		14'h2e14:	ff_dbi <= 8'h00;
		14'h2e15:	ff_dbi <= 8'h00;
		14'h2e16:	ff_dbi <= 8'h00;
		14'h2e17:	ff_dbi <= 8'h00;
		14'h2e18:	ff_dbi <= 8'h00;
		14'h2e19:	ff_dbi <= 8'h00;
		14'h2e1a:	ff_dbi <= 8'h00;
		14'h2e1b:	ff_dbi <= 8'h00;
		14'h2e1c:	ff_dbi <= 8'h00;
		14'h2e1d:	ff_dbi <= 8'h00;
		14'h2e1e:	ff_dbi <= 8'h00;
		14'h2e1f:	ff_dbi <= 8'h00;
		14'h2e20:	ff_dbi <= 8'h00;
		14'h2e21:	ff_dbi <= 8'h00;
		14'h2e22:	ff_dbi <= 8'h00;
		14'h2e23:	ff_dbi <= 8'h00;
		14'h2e24:	ff_dbi <= 8'h00;
		14'h2e25:	ff_dbi <= 8'h00;
		14'h2e26:	ff_dbi <= 8'h00;
		14'h2e27:	ff_dbi <= 8'h00;
		14'h2e28:	ff_dbi <= 8'h00;
		14'h2e29:	ff_dbi <= 8'h00;
		14'h2e2a:	ff_dbi <= 8'h00;
		14'h2e2b:	ff_dbi <= 8'h00;
		14'h2e2c:	ff_dbi <= 8'h00;
		14'h2e2d:	ff_dbi <= 8'h00;
		14'h2e2e:	ff_dbi <= 8'h00;
		14'h2e2f:	ff_dbi <= 8'h00;
		14'h2e30:	ff_dbi <= 8'h00;
		14'h2e31:	ff_dbi <= 8'h00;
		14'h2e32:	ff_dbi <= 8'h00;
		14'h2e33:	ff_dbi <= 8'h00;
		14'h2e34:	ff_dbi <= 8'h00;
		14'h2e35:	ff_dbi <= 8'h00;
		14'h2e36:	ff_dbi <= 8'h00;
		14'h2e37:	ff_dbi <= 8'h00;
		14'h2e38:	ff_dbi <= 8'h00;
		14'h2e39:	ff_dbi <= 8'h00;
		14'h2e3a:	ff_dbi <= 8'h00;
		14'h2e3b:	ff_dbi <= 8'h00;
		14'h2e3c:	ff_dbi <= 8'h00;
		14'h2e3d:	ff_dbi <= 8'h00;
		14'h2e3e:	ff_dbi <= 8'h00;
		14'h2e3f:	ff_dbi <= 8'h00;
		14'h2e40:	ff_dbi <= 8'h00;
		14'h2e41:	ff_dbi <= 8'h00;
		14'h2e42:	ff_dbi <= 8'h00;
		14'h2e43:	ff_dbi <= 8'h00;
		14'h2e44:	ff_dbi <= 8'h00;
		14'h2e45:	ff_dbi <= 8'h00;
		14'h2e46:	ff_dbi <= 8'h00;
		14'h2e47:	ff_dbi <= 8'h00;
		14'h2e48:	ff_dbi <= 8'h00;
		14'h2e49:	ff_dbi <= 8'h00;
		14'h2e4a:	ff_dbi <= 8'h00;
		14'h2e4b:	ff_dbi <= 8'h00;
		14'h2e4c:	ff_dbi <= 8'h00;
		14'h2e4d:	ff_dbi <= 8'h00;
		14'h2e4e:	ff_dbi <= 8'h00;
		14'h2e4f:	ff_dbi <= 8'h00;
		14'h2e50:	ff_dbi <= 8'h00;
		14'h2e51:	ff_dbi <= 8'h00;
		14'h2e52:	ff_dbi <= 8'h00;
		14'h2e53:	ff_dbi <= 8'h00;
		14'h2e54:	ff_dbi <= 8'h00;
		14'h2e55:	ff_dbi <= 8'h00;
		14'h2e56:	ff_dbi <= 8'h00;
		14'h2e57:	ff_dbi <= 8'h00;
		14'h2e58:	ff_dbi <= 8'h00;
		14'h2e59:	ff_dbi <= 8'h00;
		14'h2e5a:	ff_dbi <= 8'h00;
		14'h2e5b:	ff_dbi <= 8'h00;
		14'h2e5c:	ff_dbi <= 8'h00;
		14'h2e5d:	ff_dbi <= 8'h00;
		14'h2e5e:	ff_dbi <= 8'h00;
		14'h2e5f:	ff_dbi <= 8'h00;
		14'h2e60:	ff_dbi <= 8'h00;
		14'h2e61:	ff_dbi <= 8'h00;
		14'h2e62:	ff_dbi <= 8'h00;
		14'h2e63:	ff_dbi <= 8'h00;
		14'h2e64:	ff_dbi <= 8'h00;
		14'h2e65:	ff_dbi <= 8'h00;
		14'h2e66:	ff_dbi <= 8'h00;
		14'h2e67:	ff_dbi <= 8'h00;
		14'h2e68:	ff_dbi <= 8'h00;
		14'h2e69:	ff_dbi <= 8'h00;
		14'h2e6a:	ff_dbi <= 8'h00;
		14'h2e6b:	ff_dbi <= 8'h00;
		14'h2e6c:	ff_dbi <= 8'h00;
		14'h2e6d:	ff_dbi <= 8'h00;
		14'h2e6e:	ff_dbi <= 8'h00;
		14'h2e6f:	ff_dbi <= 8'h00;
		14'h2e70:	ff_dbi <= 8'h00;
		14'h2e71:	ff_dbi <= 8'h00;
		14'h2e72:	ff_dbi <= 8'h00;
		14'h2e73:	ff_dbi <= 8'h00;
		14'h2e74:	ff_dbi <= 8'h00;
		14'h2e75:	ff_dbi <= 8'h00;
		14'h2e76:	ff_dbi <= 8'h00;
		14'h2e77:	ff_dbi <= 8'h00;
		14'h2e78:	ff_dbi <= 8'h00;
		14'h2e79:	ff_dbi <= 8'h00;
		14'h2e7a:	ff_dbi <= 8'h00;
		14'h2e7b:	ff_dbi <= 8'h00;
		14'h2e7c:	ff_dbi <= 8'h00;
		14'h2e7d:	ff_dbi <= 8'h00;
		14'h2e7e:	ff_dbi <= 8'h00;
		14'h2e7f:	ff_dbi <= 8'h00;
		14'h2e80:	ff_dbi <= 8'h00;
		14'h2e81:	ff_dbi <= 8'h00;
		14'h2e82:	ff_dbi <= 8'h00;
		14'h2e83:	ff_dbi <= 8'h00;
		14'h2e84:	ff_dbi <= 8'h00;
		14'h2e85:	ff_dbi <= 8'h00;
		14'h2e86:	ff_dbi <= 8'h00;
		14'h2e87:	ff_dbi <= 8'h00;
		14'h2e88:	ff_dbi <= 8'h00;
		14'h2e89:	ff_dbi <= 8'h00;
		14'h2e8a:	ff_dbi <= 8'h00;
		14'h2e8b:	ff_dbi <= 8'h00;
		14'h2e8c:	ff_dbi <= 8'h00;
		14'h2e8d:	ff_dbi <= 8'h00;
		14'h2e8e:	ff_dbi <= 8'h00;
		14'h2e8f:	ff_dbi <= 8'h00;
		14'h2e90:	ff_dbi <= 8'h00;
		14'h2e91:	ff_dbi <= 8'h00;
		14'h2e92:	ff_dbi <= 8'h00;
		14'h2e93:	ff_dbi <= 8'h00;
		14'h2e94:	ff_dbi <= 8'h00;
		14'h2e95:	ff_dbi <= 8'h00;
		14'h2e96:	ff_dbi <= 8'h00;
		14'h2e97:	ff_dbi <= 8'h00;
		14'h2e98:	ff_dbi <= 8'h00;
		14'h2e99:	ff_dbi <= 8'h00;
		14'h2e9a:	ff_dbi <= 8'h00;
		14'h2e9b:	ff_dbi <= 8'h00;
		14'h2e9c:	ff_dbi <= 8'h00;
		14'h2e9d:	ff_dbi <= 8'h00;
		14'h2e9e:	ff_dbi <= 8'h00;
		14'h2e9f:	ff_dbi <= 8'h00;
		14'h2ea0:	ff_dbi <= 8'h00;
		14'h2ea1:	ff_dbi <= 8'h00;
		14'h2ea2:	ff_dbi <= 8'h00;
		14'h2ea3:	ff_dbi <= 8'h00;
		14'h2ea4:	ff_dbi <= 8'h00;
		14'h2ea5:	ff_dbi <= 8'h00;
		14'h2ea6:	ff_dbi <= 8'h00;
		14'h2ea7:	ff_dbi <= 8'h00;
		14'h2ea8:	ff_dbi <= 8'h00;
		14'h2ea9:	ff_dbi <= 8'h00;
		14'h2eaa:	ff_dbi <= 8'h00;
		14'h2eab:	ff_dbi <= 8'h00;
		14'h2eac:	ff_dbi <= 8'h00;
		14'h2ead:	ff_dbi <= 8'h00;
		14'h2eae:	ff_dbi <= 8'h00;
		14'h2eaf:	ff_dbi <= 8'h00;
		14'h2eb0:	ff_dbi <= 8'h00;
		14'h2eb1:	ff_dbi <= 8'h00;
		14'h2eb2:	ff_dbi <= 8'h00;
		14'h2eb3:	ff_dbi <= 8'h00;
		14'h2eb4:	ff_dbi <= 8'h00;
		14'h2eb5:	ff_dbi <= 8'h00;
		14'h2eb6:	ff_dbi <= 8'h00;
		14'h2eb7:	ff_dbi <= 8'h00;
		14'h2eb8:	ff_dbi <= 8'h00;
		14'h2eb9:	ff_dbi <= 8'h00;
		14'h2eba:	ff_dbi <= 8'h00;
		14'h2ebb:	ff_dbi <= 8'h00;
		14'h2ebc:	ff_dbi <= 8'h00;
		14'h2ebd:	ff_dbi <= 8'h00;
		14'h2ebe:	ff_dbi <= 8'h00;
		14'h2ebf:	ff_dbi <= 8'h00;
		14'h2ec0:	ff_dbi <= 8'h00;
		14'h2ec1:	ff_dbi <= 8'h00;
		14'h2ec2:	ff_dbi <= 8'h00;
		14'h2ec3:	ff_dbi <= 8'h00;
		14'h2ec4:	ff_dbi <= 8'h00;
		14'h2ec5:	ff_dbi <= 8'h00;
		14'h2ec6:	ff_dbi <= 8'h00;
		14'h2ec7:	ff_dbi <= 8'h00;
		14'h2ec8:	ff_dbi <= 8'h00;
		14'h2ec9:	ff_dbi <= 8'h00;
		14'h2eca:	ff_dbi <= 8'h00;
		14'h2ecb:	ff_dbi <= 8'h00;
		14'h2ecc:	ff_dbi <= 8'h00;
		14'h2ecd:	ff_dbi <= 8'h00;
		14'h2ece:	ff_dbi <= 8'h00;
		14'h2ecf:	ff_dbi <= 8'h00;
		14'h2ed0:	ff_dbi <= 8'h00;
		14'h2ed1:	ff_dbi <= 8'h00;
		14'h2ed2:	ff_dbi <= 8'h00;
		14'h2ed3:	ff_dbi <= 8'h00;
		14'h2ed4:	ff_dbi <= 8'h00;
		14'h2ed5:	ff_dbi <= 8'h00;
		14'h2ed6:	ff_dbi <= 8'h00;
		14'h2ed7:	ff_dbi <= 8'h00;
		14'h2ed8:	ff_dbi <= 8'h00;
		14'h2ed9:	ff_dbi <= 8'h00;
		14'h2eda:	ff_dbi <= 8'h00;
		14'h2edb:	ff_dbi <= 8'h00;
		14'h2edc:	ff_dbi <= 8'h00;
		14'h2edd:	ff_dbi <= 8'h00;
		14'h2ede:	ff_dbi <= 8'h00;
		14'h2edf:	ff_dbi <= 8'h00;
		14'h2ee0:	ff_dbi <= 8'h00;
		14'h2ee1:	ff_dbi <= 8'h00;
		14'h2ee2:	ff_dbi <= 8'h00;
		14'h2ee3:	ff_dbi <= 8'h00;
		14'h2ee4:	ff_dbi <= 8'h00;
		14'h2ee5:	ff_dbi <= 8'h00;
		14'h2ee6:	ff_dbi <= 8'h00;
		14'h2ee7:	ff_dbi <= 8'h00;
		14'h2ee8:	ff_dbi <= 8'h00;
		14'h2ee9:	ff_dbi <= 8'h00;
		14'h2eea:	ff_dbi <= 8'h00;
		14'h2eeb:	ff_dbi <= 8'h00;
		14'h2eec:	ff_dbi <= 8'h00;
		14'h2eed:	ff_dbi <= 8'h00;
		14'h2eee:	ff_dbi <= 8'h00;
		14'h2eef:	ff_dbi <= 8'h00;
		14'h2ef0:	ff_dbi <= 8'h00;
		14'h2ef1:	ff_dbi <= 8'h00;
		14'h2ef2:	ff_dbi <= 8'h00;
		14'h2ef3:	ff_dbi <= 8'h00;
		14'h2ef4:	ff_dbi <= 8'h00;
		14'h2ef5:	ff_dbi <= 8'h00;
		14'h2ef6:	ff_dbi <= 8'h00;
		14'h2ef7:	ff_dbi <= 8'h00;
		14'h2ef8:	ff_dbi <= 8'h00;
		14'h2ef9:	ff_dbi <= 8'h00;
		14'h2efa:	ff_dbi <= 8'h00;
		14'h2efb:	ff_dbi <= 8'h00;
		14'h2efc:	ff_dbi <= 8'h00;
		14'h2efd:	ff_dbi <= 8'h00;
		14'h2efe:	ff_dbi <= 8'h00;
		14'h2eff:	ff_dbi <= 8'h00;
		14'h2f00:	ff_dbi <= 8'h00;
		14'h2f01:	ff_dbi <= 8'h00;
		14'h2f02:	ff_dbi <= 8'h00;
		14'h2f03:	ff_dbi <= 8'h00;
		14'h2f04:	ff_dbi <= 8'h00;
		14'h2f05:	ff_dbi <= 8'h00;
		14'h2f06:	ff_dbi <= 8'h00;
		14'h2f07:	ff_dbi <= 8'h00;
		14'h2f08:	ff_dbi <= 8'h00;
		14'h2f09:	ff_dbi <= 8'h00;
		14'h2f0a:	ff_dbi <= 8'h00;
		14'h2f0b:	ff_dbi <= 8'h00;
		14'h2f0c:	ff_dbi <= 8'h00;
		14'h2f0d:	ff_dbi <= 8'h00;
		14'h2f0e:	ff_dbi <= 8'h00;
		14'h2f0f:	ff_dbi <= 8'h00;
		14'h2f10:	ff_dbi <= 8'h00;
		14'h2f11:	ff_dbi <= 8'h00;
		14'h2f12:	ff_dbi <= 8'h00;
		14'h2f13:	ff_dbi <= 8'h00;
		14'h2f14:	ff_dbi <= 8'h00;
		14'h2f15:	ff_dbi <= 8'h00;
		14'h2f16:	ff_dbi <= 8'h00;
		14'h2f17:	ff_dbi <= 8'h00;
		14'h2f18:	ff_dbi <= 8'h00;
		14'h2f19:	ff_dbi <= 8'h00;
		14'h2f1a:	ff_dbi <= 8'h00;
		14'h2f1b:	ff_dbi <= 8'h00;
		14'h2f1c:	ff_dbi <= 8'h00;
		14'h2f1d:	ff_dbi <= 8'h00;
		14'h2f1e:	ff_dbi <= 8'h00;
		14'h2f1f:	ff_dbi <= 8'h00;
		14'h2f20:	ff_dbi <= 8'h00;
		14'h2f21:	ff_dbi <= 8'h00;
		14'h2f22:	ff_dbi <= 8'h00;
		14'h2f23:	ff_dbi <= 8'h00;
		14'h2f24:	ff_dbi <= 8'h00;
		14'h2f25:	ff_dbi <= 8'h00;
		14'h2f26:	ff_dbi <= 8'h00;
		14'h2f27:	ff_dbi <= 8'h00;
		14'h2f28:	ff_dbi <= 8'h00;
		14'h2f29:	ff_dbi <= 8'h00;
		14'h2f2a:	ff_dbi <= 8'h00;
		14'h2f2b:	ff_dbi <= 8'h00;
		14'h2f2c:	ff_dbi <= 8'h00;
		14'h2f2d:	ff_dbi <= 8'h00;
		14'h2f2e:	ff_dbi <= 8'h00;
		14'h2f2f:	ff_dbi <= 8'h00;
		14'h2f30:	ff_dbi <= 8'h00;
		14'h2f31:	ff_dbi <= 8'h00;
		14'h2f32:	ff_dbi <= 8'h00;
		14'h2f33:	ff_dbi <= 8'h00;
		14'h2f34:	ff_dbi <= 8'h00;
		14'h2f35:	ff_dbi <= 8'h00;
		14'h2f36:	ff_dbi <= 8'h00;
		14'h2f37:	ff_dbi <= 8'h00;
		14'h2f38:	ff_dbi <= 8'h00;
		14'h2f39:	ff_dbi <= 8'h00;
		14'h2f3a:	ff_dbi <= 8'h00;
		14'h2f3b:	ff_dbi <= 8'h00;
		14'h2f3c:	ff_dbi <= 8'h00;
		14'h2f3d:	ff_dbi <= 8'h00;
		14'h2f3e:	ff_dbi <= 8'h00;
		14'h2f3f:	ff_dbi <= 8'h00;
		14'h2f40:	ff_dbi <= 8'h00;
		14'h2f41:	ff_dbi <= 8'h00;
		14'h2f42:	ff_dbi <= 8'h00;
		14'h2f43:	ff_dbi <= 8'h00;
		14'h2f44:	ff_dbi <= 8'h00;
		14'h2f45:	ff_dbi <= 8'h00;
		14'h2f46:	ff_dbi <= 8'h00;
		14'h2f47:	ff_dbi <= 8'h00;
		14'h2f48:	ff_dbi <= 8'h00;
		14'h2f49:	ff_dbi <= 8'h00;
		14'h2f4a:	ff_dbi <= 8'h00;
		14'h2f4b:	ff_dbi <= 8'h00;
		14'h2f4c:	ff_dbi <= 8'h00;
		14'h2f4d:	ff_dbi <= 8'h00;
		14'h2f4e:	ff_dbi <= 8'h00;
		14'h2f4f:	ff_dbi <= 8'h00;
		14'h2f50:	ff_dbi <= 8'h00;
		14'h2f51:	ff_dbi <= 8'h00;
		14'h2f52:	ff_dbi <= 8'h00;
		14'h2f53:	ff_dbi <= 8'h00;
		14'h2f54:	ff_dbi <= 8'h00;
		14'h2f55:	ff_dbi <= 8'h00;
		14'h2f56:	ff_dbi <= 8'h00;
		14'h2f57:	ff_dbi <= 8'h00;
		14'h2f58:	ff_dbi <= 8'h00;
		14'h2f59:	ff_dbi <= 8'h00;
		14'h2f5a:	ff_dbi <= 8'h00;
		14'h2f5b:	ff_dbi <= 8'h00;
		14'h2f5c:	ff_dbi <= 8'h00;
		14'h2f5d:	ff_dbi <= 8'h00;
		14'h2f5e:	ff_dbi <= 8'h00;
		14'h2f5f:	ff_dbi <= 8'h00;
		14'h2f60:	ff_dbi <= 8'h00;
		14'h2f61:	ff_dbi <= 8'h00;
		14'h2f62:	ff_dbi <= 8'h00;
		14'h2f63:	ff_dbi <= 8'h00;
		14'h2f64:	ff_dbi <= 8'h00;
		14'h2f65:	ff_dbi <= 8'h00;
		14'h2f66:	ff_dbi <= 8'h00;
		14'h2f67:	ff_dbi <= 8'h00;
		14'h2f68:	ff_dbi <= 8'h00;
		14'h2f69:	ff_dbi <= 8'h00;
		14'h2f6a:	ff_dbi <= 8'h00;
		14'h2f6b:	ff_dbi <= 8'h00;
		14'h2f6c:	ff_dbi <= 8'h00;
		14'h2f6d:	ff_dbi <= 8'h00;
		14'h2f6e:	ff_dbi <= 8'h00;
		14'h2f6f:	ff_dbi <= 8'h00;
		14'h2f70:	ff_dbi <= 8'h00;
		14'h2f71:	ff_dbi <= 8'h00;
		14'h2f72:	ff_dbi <= 8'h00;
		14'h2f73:	ff_dbi <= 8'h00;
		14'h2f74:	ff_dbi <= 8'h00;
		14'h2f75:	ff_dbi <= 8'h00;
		14'h2f76:	ff_dbi <= 8'h00;
		14'h2f77:	ff_dbi <= 8'h00;
		14'h2f78:	ff_dbi <= 8'h00;
		14'h2f79:	ff_dbi <= 8'h00;
		14'h2f7a:	ff_dbi <= 8'h00;
		14'h2f7b:	ff_dbi <= 8'h00;
		14'h2f7c:	ff_dbi <= 8'h00;
		14'h2f7d:	ff_dbi <= 8'h00;
		14'h2f7e:	ff_dbi <= 8'h00;
		14'h2f7f:	ff_dbi <= 8'h00;
		14'h2f80:	ff_dbi <= 8'h00;
		14'h2f81:	ff_dbi <= 8'h00;
		14'h2f82:	ff_dbi <= 8'h00;
		14'h2f83:	ff_dbi <= 8'h00;
		14'h2f84:	ff_dbi <= 8'h00;
		14'h2f85:	ff_dbi <= 8'h00;
		14'h2f86:	ff_dbi <= 8'h00;
		14'h2f87:	ff_dbi <= 8'h00;
		14'h2f88:	ff_dbi <= 8'h00;
		14'h2f89:	ff_dbi <= 8'h00;
		14'h2f8a:	ff_dbi <= 8'h00;
		14'h2f8b:	ff_dbi <= 8'h00;
		14'h2f8c:	ff_dbi <= 8'h00;
		14'h2f8d:	ff_dbi <= 8'h00;
		14'h2f8e:	ff_dbi <= 8'h00;
		14'h2f8f:	ff_dbi <= 8'h00;
		14'h2f90:	ff_dbi <= 8'h00;
		14'h2f91:	ff_dbi <= 8'h00;
		14'h2f92:	ff_dbi <= 8'h00;
		14'h2f93:	ff_dbi <= 8'h00;
		14'h2f94:	ff_dbi <= 8'h00;
		14'h2f95:	ff_dbi <= 8'h00;
		14'h2f96:	ff_dbi <= 8'h00;
		14'h2f97:	ff_dbi <= 8'h00;
		14'h2f98:	ff_dbi <= 8'h00;
		14'h2f99:	ff_dbi <= 8'h00;
		14'h2f9a:	ff_dbi <= 8'h00;
		14'h2f9b:	ff_dbi <= 8'h00;
		14'h2f9c:	ff_dbi <= 8'h00;
		14'h2f9d:	ff_dbi <= 8'h00;
		14'h2f9e:	ff_dbi <= 8'h00;
		14'h2f9f:	ff_dbi <= 8'h00;
		14'h2fa0:	ff_dbi <= 8'h00;
		14'h2fa1:	ff_dbi <= 8'h00;
		14'h2fa2:	ff_dbi <= 8'h00;
		14'h2fa3:	ff_dbi <= 8'h00;
		14'h2fa4:	ff_dbi <= 8'h00;
		14'h2fa5:	ff_dbi <= 8'h00;
		14'h2fa6:	ff_dbi <= 8'h00;
		14'h2fa7:	ff_dbi <= 8'h00;
		14'h2fa8:	ff_dbi <= 8'h00;
		14'h2fa9:	ff_dbi <= 8'h00;
		14'h2faa:	ff_dbi <= 8'h00;
		14'h2fab:	ff_dbi <= 8'h00;
		14'h2fac:	ff_dbi <= 8'h00;
		14'h2fad:	ff_dbi <= 8'h00;
		14'h2fae:	ff_dbi <= 8'h00;
		14'h2faf:	ff_dbi <= 8'h00;
		14'h2fb0:	ff_dbi <= 8'h00;
		14'h2fb1:	ff_dbi <= 8'h00;
		14'h2fb2:	ff_dbi <= 8'h00;
		14'h2fb3:	ff_dbi <= 8'h00;
		14'h2fb4:	ff_dbi <= 8'h00;
		14'h2fb5:	ff_dbi <= 8'h00;
		14'h2fb6:	ff_dbi <= 8'h00;
		14'h2fb7:	ff_dbi <= 8'h00;
		14'h2fb8:	ff_dbi <= 8'h00;
		14'h2fb9:	ff_dbi <= 8'h00;
		14'h2fba:	ff_dbi <= 8'h00;
		14'h2fbb:	ff_dbi <= 8'h00;
		14'h2fbc:	ff_dbi <= 8'h00;
		14'h2fbd:	ff_dbi <= 8'h00;
		14'h2fbe:	ff_dbi <= 8'h00;
		14'h2fbf:	ff_dbi <= 8'h00;
		14'h2fc0:	ff_dbi <= 8'h00;
		14'h2fc1:	ff_dbi <= 8'h00;
		14'h2fc2:	ff_dbi <= 8'h00;
		14'h2fc3:	ff_dbi <= 8'h00;
		14'h2fc4:	ff_dbi <= 8'h00;
		14'h2fc5:	ff_dbi <= 8'h00;
		14'h2fc6:	ff_dbi <= 8'h00;
		14'h2fc7:	ff_dbi <= 8'h00;
		14'h2fc8:	ff_dbi <= 8'h00;
		14'h2fc9:	ff_dbi <= 8'h00;
		14'h2fca:	ff_dbi <= 8'h00;
		14'h2fcb:	ff_dbi <= 8'h00;
		14'h2fcc:	ff_dbi <= 8'h00;
		14'h2fcd:	ff_dbi <= 8'h00;
		14'h2fce:	ff_dbi <= 8'h00;
		14'h2fcf:	ff_dbi <= 8'h00;
		14'h2fd0:	ff_dbi <= 8'h00;
		14'h2fd1:	ff_dbi <= 8'h00;
		14'h2fd2:	ff_dbi <= 8'h00;
		14'h2fd3:	ff_dbi <= 8'h00;
		14'h2fd4:	ff_dbi <= 8'h00;
		14'h2fd5:	ff_dbi <= 8'h00;
		14'h2fd6:	ff_dbi <= 8'h00;
		14'h2fd7:	ff_dbi <= 8'h00;
		14'h2fd8:	ff_dbi <= 8'h00;
		14'h2fd9:	ff_dbi <= 8'h00;
		14'h2fda:	ff_dbi <= 8'h00;
		14'h2fdb:	ff_dbi <= 8'h00;
		14'h2fdc:	ff_dbi <= 8'h00;
		14'h2fdd:	ff_dbi <= 8'h00;
		14'h2fde:	ff_dbi <= 8'h00;
		14'h2fdf:	ff_dbi <= 8'h00;
		14'h2fe0:	ff_dbi <= 8'h00;
		14'h2fe1:	ff_dbi <= 8'h00;
		14'h2fe2:	ff_dbi <= 8'h00;
		14'h2fe3:	ff_dbi <= 8'h00;
		14'h2fe4:	ff_dbi <= 8'h00;
		14'h2fe5:	ff_dbi <= 8'h00;
		14'h2fe6:	ff_dbi <= 8'h00;
		14'h2fe7:	ff_dbi <= 8'h00;
		14'h2fe8:	ff_dbi <= 8'h00;
		14'h2fe9:	ff_dbi <= 8'h00;
		14'h2fea:	ff_dbi <= 8'h00;
		14'h2feb:	ff_dbi <= 8'h00;
		14'h2fec:	ff_dbi <= 8'h00;
		14'h2fed:	ff_dbi <= 8'h00;
		14'h2fee:	ff_dbi <= 8'h00;
		14'h2fef:	ff_dbi <= 8'h00;
		14'h2ff0:	ff_dbi <= 8'h00;
		14'h2ff1:	ff_dbi <= 8'h00;
		14'h2ff2:	ff_dbi <= 8'h00;
		14'h2ff3:	ff_dbi <= 8'h00;
		14'h2ff4:	ff_dbi <= 8'h00;
		14'h2ff5:	ff_dbi <= 8'h00;
		14'h2ff6:	ff_dbi <= 8'h00;
		14'h2ff7:	ff_dbi <= 8'h00;
		14'h2ff8:	ff_dbi <= 8'h00;
		14'h2ff9:	ff_dbi <= 8'h00;
		14'h2ffa:	ff_dbi <= 8'h00;
		14'h2ffb:	ff_dbi <= 8'h00;
		14'h2ffc:	ff_dbi <= 8'h00;
		14'h2ffd:	ff_dbi <= 8'h00;
		14'h2ffe:	ff_dbi <= 8'h00;
		14'h2fff:	ff_dbi <= 8'h00;
		14'h3000:	ff_dbi <= 8'h00;
		14'h3001:	ff_dbi <= 8'h00;
		14'h3002:	ff_dbi <= 8'h00;
		14'h3003:	ff_dbi <= 8'h00;
		14'h3004:	ff_dbi <= 8'h00;
		14'h3005:	ff_dbi <= 8'h00;
		14'h3006:	ff_dbi <= 8'h00;
		14'h3007:	ff_dbi <= 8'h00;
		14'h3008:	ff_dbi <= 8'h00;
		14'h3009:	ff_dbi <= 8'h00;
		14'h300a:	ff_dbi <= 8'h00;
		14'h300b:	ff_dbi <= 8'h00;
		14'h300c:	ff_dbi <= 8'h00;
		14'h300d:	ff_dbi <= 8'h00;
		14'h300e:	ff_dbi <= 8'h00;
		14'h300f:	ff_dbi <= 8'h00;
		14'h3010:	ff_dbi <= 8'h00;
		14'h3011:	ff_dbi <= 8'h00;
		14'h3012:	ff_dbi <= 8'h00;
		14'h3013:	ff_dbi <= 8'h00;
		14'h3014:	ff_dbi <= 8'h00;
		14'h3015:	ff_dbi <= 8'h00;
		14'h3016:	ff_dbi <= 8'h00;
		14'h3017:	ff_dbi <= 8'h00;
		14'h3018:	ff_dbi <= 8'h00;
		14'h3019:	ff_dbi <= 8'h00;
		14'h301a:	ff_dbi <= 8'h00;
		14'h301b:	ff_dbi <= 8'h00;
		14'h301c:	ff_dbi <= 8'h00;
		14'h301d:	ff_dbi <= 8'h00;
		14'h301e:	ff_dbi <= 8'h00;
		14'h301f:	ff_dbi <= 8'h00;
		14'h3020:	ff_dbi <= 8'h00;
		14'h3021:	ff_dbi <= 8'h00;
		14'h3022:	ff_dbi <= 8'h00;
		14'h3023:	ff_dbi <= 8'h00;
		14'h3024:	ff_dbi <= 8'h00;
		14'h3025:	ff_dbi <= 8'h00;
		14'h3026:	ff_dbi <= 8'h00;
		14'h3027:	ff_dbi <= 8'h00;
		14'h3028:	ff_dbi <= 8'h00;
		14'h3029:	ff_dbi <= 8'h00;
		14'h302a:	ff_dbi <= 8'h00;
		14'h302b:	ff_dbi <= 8'h00;
		14'h302c:	ff_dbi <= 8'h00;
		14'h302d:	ff_dbi <= 8'h00;
		14'h302e:	ff_dbi <= 8'h00;
		14'h302f:	ff_dbi <= 8'h00;
		14'h3030:	ff_dbi <= 8'h00;
		14'h3031:	ff_dbi <= 8'h00;
		14'h3032:	ff_dbi <= 8'h00;
		14'h3033:	ff_dbi <= 8'h00;
		14'h3034:	ff_dbi <= 8'h00;
		14'h3035:	ff_dbi <= 8'h00;
		14'h3036:	ff_dbi <= 8'h00;
		14'h3037:	ff_dbi <= 8'h00;
		14'h3038:	ff_dbi <= 8'h00;
		14'h3039:	ff_dbi <= 8'h00;
		14'h303a:	ff_dbi <= 8'h00;
		14'h303b:	ff_dbi <= 8'h00;
		14'h303c:	ff_dbi <= 8'h00;
		14'h303d:	ff_dbi <= 8'h00;
		14'h303e:	ff_dbi <= 8'h00;
		14'h303f:	ff_dbi <= 8'h00;
		14'h3040:	ff_dbi <= 8'h00;
		14'h3041:	ff_dbi <= 8'h00;
		14'h3042:	ff_dbi <= 8'h00;
		14'h3043:	ff_dbi <= 8'h00;
		14'h3044:	ff_dbi <= 8'h00;
		14'h3045:	ff_dbi <= 8'h00;
		14'h3046:	ff_dbi <= 8'h00;
		14'h3047:	ff_dbi <= 8'h00;
		14'h3048:	ff_dbi <= 8'h00;
		14'h3049:	ff_dbi <= 8'h00;
		14'h304a:	ff_dbi <= 8'h00;
		14'h304b:	ff_dbi <= 8'h00;
		14'h304c:	ff_dbi <= 8'h00;
		14'h304d:	ff_dbi <= 8'h00;
		14'h304e:	ff_dbi <= 8'h00;
		14'h304f:	ff_dbi <= 8'h00;
		14'h3050:	ff_dbi <= 8'h00;
		14'h3051:	ff_dbi <= 8'h00;
		14'h3052:	ff_dbi <= 8'h00;
		14'h3053:	ff_dbi <= 8'h00;
		14'h3054:	ff_dbi <= 8'h00;
		14'h3055:	ff_dbi <= 8'h00;
		14'h3056:	ff_dbi <= 8'h00;
		14'h3057:	ff_dbi <= 8'h00;
		14'h3058:	ff_dbi <= 8'h00;
		14'h3059:	ff_dbi <= 8'h00;
		14'h305a:	ff_dbi <= 8'h00;
		14'h305b:	ff_dbi <= 8'h00;
		14'h305c:	ff_dbi <= 8'h00;
		14'h305d:	ff_dbi <= 8'h00;
		14'h305e:	ff_dbi <= 8'h00;
		14'h305f:	ff_dbi <= 8'h00;
		14'h3060:	ff_dbi <= 8'h00;
		14'h3061:	ff_dbi <= 8'h00;
		14'h3062:	ff_dbi <= 8'h00;
		14'h3063:	ff_dbi <= 8'h00;
		14'h3064:	ff_dbi <= 8'h00;
		14'h3065:	ff_dbi <= 8'h00;
		14'h3066:	ff_dbi <= 8'h00;
		14'h3067:	ff_dbi <= 8'h00;
		14'h3068:	ff_dbi <= 8'h00;
		14'h3069:	ff_dbi <= 8'h00;
		14'h306a:	ff_dbi <= 8'h00;
		14'h306b:	ff_dbi <= 8'h00;
		14'h306c:	ff_dbi <= 8'h00;
		14'h306d:	ff_dbi <= 8'h00;
		14'h306e:	ff_dbi <= 8'h00;
		14'h306f:	ff_dbi <= 8'h00;
		14'h3070:	ff_dbi <= 8'h00;
		14'h3071:	ff_dbi <= 8'h00;
		14'h3072:	ff_dbi <= 8'h00;
		14'h3073:	ff_dbi <= 8'h00;
		14'h3074:	ff_dbi <= 8'h00;
		14'h3075:	ff_dbi <= 8'h00;
		14'h3076:	ff_dbi <= 8'h00;
		14'h3077:	ff_dbi <= 8'h00;
		14'h3078:	ff_dbi <= 8'h00;
		14'h3079:	ff_dbi <= 8'h00;
		14'h307a:	ff_dbi <= 8'h00;
		14'h307b:	ff_dbi <= 8'h00;
		14'h307c:	ff_dbi <= 8'h00;
		14'h307d:	ff_dbi <= 8'h00;
		14'h307e:	ff_dbi <= 8'h00;
		14'h307f:	ff_dbi <= 8'h00;
		14'h3080:	ff_dbi <= 8'h00;
		14'h3081:	ff_dbi <= 8'h00;
		14'h3082:	ff_dbi <= 8'h00;
		14'h3083:	ff_dbi <= 8'h00;
		14'h3084:	ff_dbi <= 8'h00;
		14'h3085:	ff_dbi <= 8'h00;
		14'h3086:	ff_dbi <= 8'h00;
		14'h3087:	ff_dbi <= 8'h00;
		14'h3088:	ff_dbi <= 8'h00;
		14'h3089:	ff_dbi <= 8'h00;
		14'h308a:	ff_dbi <= 8'h00;
		14'h308b:	ff_dbi <= 8'h00;
		14'h308c:	ff_dbi <= 8'h00;
		14'h308d:	ff_dbi <= 8'h00;
		14'h308e:	ff_dbi <= 8'h00;
		14'h308f:	ff_dbi <= 8'h00;
		14'h3090:	ff_dbi <= 8'h00;
		14'h3091:	ff_dbi <= 8'h00;
		14'h3092:	ff_dbi <= 8'h00;
		14'h3093:	ff_dbi <= 8'h00;
		14'h3094:	ff_dbi <= 8'h00;
		14'h3095:	ff_dbi <= 8'h00;
		14'h3096:	ff_dbi <= 8'h00;
		14'h3097:	ff_dbi <= 8'h00;
		14'h3098:	ff_dbi <= 8'h00;
		14'h3099:	ff_dbi <= 8'h00;
		14'h309a:	ff_dbi <= 8'h00;
		14'h309b:	ff_dbi <= 8'h00;
		14'h309c:	ff_dbi <= 8'h00;
		14'h309d:	ff_dbi <= 8'h00;
		14'h309e:	ff_dbi <= 8'h00;
		14'h309f:	ff_dbi <= 8'h00;
		14'h30a0:	ff_dbi <= 8'h00;
		14'h30a1:	ff_dbi <= 8'h00;
		14'h30a2:	ff_dbi <= 8'h00;
		14'h30a3:	ff_dbi <= 8'h00;
		14'h30a4:	ff_dbi <= 8'h00;
		14'h30a5:	ff_dbi <= 8'h00;
		14'h30a6:	ff_dbi <= 8'h00;
		14'h30a7:	ff_dbi <= 8'h00;
		14'h30a8:	ff_dbi <= 8'h00;
		14'h30a9:	ff_dbi <= 8'h00;
		14'h30aa:	ff_dbi <= 8'h00;
		14'h30ab:	ff_dbi <= 8'h00;
		14'h30ac:	ff_dbi <= 8'h00;
		14'h30ad:	ff_dbi <= 8'h00;
		14'h30ae:	ff_dbi <= 8'h00;
		14'h30af:	ff_dbi <= 8'h00;
		14'h30b0:	ff_dbi <= 8'h00;
		14'h30b1:	ff_dbi <= 8'h00;
		14'h30b2:	ff_dbi <= 8'h00;
		14'h30b3:	ff_dbi <= 8'h00;
		14'h30b4:	ff_dbi <= 8'h00;
		14'h30b5:	ff_dbi <= 8'h00;
		14'h30b6:	ff_dbi <= 8'h00;
		14'h30b7:	ff_dbi <= 8'h00;
		14'h30b8:	ff_dbi <= 8'h00;
		14'h30b9:	ff_dbi <= 8'h00;
		14'h30ba:	ff_dbi <= 8'h00;
		14'h30bb:	ff_dbi <= 8'h00;
		14'h30bc:	ff_dbi <= 8'h00;
		14'h30bd:	ff_dbi <= 8'h00;
		14'h30be:	ff_dbi <= 8'h00;
		14'h30bf:	ff_dbi <= 8'h00;
		14'h30c0:	ff_dbi <= 8'h00;
		14'h30c1:	ff_dbi <= 8'h00;
		14'h30c2:	ff_dbi <= 8'h00;
		14'h30c3:	ff_dbi <= 8'h00;
		14'h30c4:	ff_dbi <= 8'h00;
		14'h30c5:	ff_dbi <= 8'h00;
		14'h30c6:	ff_dbi <= 8'h00;
		14'h30c7:	ff_dbi <= 8'h00;
		14'h30c8:	ff_dbi <= 8'h00;
		14'h30c9:	ff_dbi <= 8'h00;
		14'h30ca:	ff_dbi <= 8'h00;
		14'h30cb:	ff_dbi <= 8'h00;
		14'h30cc:	ff_dbi <= 8'h00;
		14'h30cd:	ff_dbi <= 8'h00;
		14'h30ce:	ff_dbi <= 8'h00;
		14'h30cf:	ff_dbi <= 8'h00;
		14'h30d0:	ff_dbi <= 8'h00;
		14'h30d1:	ff_dbi <= 8'h00;
		14'h30d2:	ff_dbi <= 8'h00;
		14'h30d3:	ff_dbi <= 8'h00;
		14'h30d4:	ff_dbi <= 8'h00;
		14'h30d5:	ff_dbi <= 8'h00;
		14'h30d6:	ff_dbi <= 8'h00;
		14'h30d7:	ff_dbi <= 8'h00;
		14'h30d8:	ff_dbi <= 8'h00;
		14'h30d9:	ff_dbi <= 8'h00;
		14'h30da:	ff_dbi <= 8'h00;
		14'h30db:	ff_dbi <= 8'h00;
		14'h30dc:	ff_dbi <= 8'h00;
		14'h30dd:	ff_dbi <= 8'h00;
		14'h30de:	ff_dbi <= 8'h00;
		14'h30df:	ff_dbi <= 8'h00;
		14'h30e0:	ff_dbi <= 8'h00;
		14'h30e1:	ff_dbi <= 8'h00;
		14'h30e2:	ff_dbi <= 8'h00;
		14'h30e3:	ff_dbi <= 8'h00;
		14'h30e4:	ff_dbi <= 8'h00;
		14'h30e5:	ff_dbi <= 8'h00;
		14'h30e6:	ff_dbi <= 8'h00;
		14'h30e7:	ff_dbi <= 8'h00;
		14'h30e8:	ff_dbi <= 8'h00;
		14'h30e9:	ff_dbi <= 8'h00;
		14'h30ea:	ff_dbi <= 8'h00;
		14'h30eb:	ff_dbi <= 8'h00;
		14'h30ec:	ff_dbi <= 8'h00;
		14'h30ed:	ff_dbi <= 8'h00;
		14'h30ee:	ff_dbi <= 8'h00;
		14'h30ef:	ff_dbi <= 8'h00;
		14'h30f0:	ff_dbi <= 8'h00;
		14'h30f1:	ff_dbi <= 8'h00;
		14'h30f2:	ff_dbi <= 8'h00;
		14'h30f3:	ff_dbi <= 8'h00;
		14'h30f4:	ff_dbi <= 8'h00;
		14'h30f5:	ff_dbi <= 8'h00;
		14'h30f6:	ff_dbi <= 8'h00;
		14'h30f7:	ff_dbi <= 8'h00;
		14'h30f8:	ff_dbi <= 8'h00;
		14'h30f9:	ff_dbi <= 8'h00;
		14'h30fa:	ff_dbi <= 8'h00;
		14'h30fb:	ff_dbi <= 8'h00;
		14'h30fc:	ff_dbi <= 8'h00;
		14'h30fd:	ff_dbi <= 8'h00;
		14'h30fe:	ff_dbi <= 8'h00;
		14'h30ff:	ff_dbi <= 8'h00;
		14'h3100:	ff_dbi <= 8'h00;
		14'h3101:	ff_dbi <= 8'h00;
		14'h3102:	ff_dbi <= 8'h00;
		14'h3103:	ff_dbi <= 8'h00;
		14'h3104:	ff_dbi <= 8'h00;
		14'h3105:	ff_dbi <= 8'h00;
		14'h3106:	ff_dbi <= 8'h00;
		14'h3107:	ff_dbi <= 8'h00;
		14'h3108:	ff_dbi <= 8'h00;
		14'h3109:	ff_dbi <= 8'h00;
		14'h310a:	ff_dbi <= 8'h00;
		14'h310b:	ff_dbi <= 8'h00;
		14'h310c:	ff_dbi <= 8'h00;
		14'h310d:	ff_dbi <= 8'h00;
		14'h310e:	ff_dbi <= 8'h00;
		14'h310f:	ff_dbi <= 8'h00;
		14'h3110:	ff_dbi <= 8'h00;
		14'h3111:	ff_dbi <= 8'h00;
		14'h3112:	ff_dbi <= 8'h00;
		14'h3113:	ff_dbi <= 8'h00;
		14'h3114:	ff_dbi <= 8'h00;
		14'h3115:	ff_dbi <= 8'h00;
		14'h3116:	ff_dbi <= 8'h00;
		14'h3117:	ff_dbi <= 8'h00;
		14'h3118:	ff_dbi <= 8'h00;
		14'h3119:	ff_dbi <= 8'h00;
		14'h311a:	ff_dbi <= 8'h00;
		14'h311b:	ff_dbi <= 8'h00;
		14'h311c:	ff_dbi <= 8'h00;
		14'h311d:	ff_dbi <= 8'h00;
		14'h311e:	ff_dbi <= 8'h00;
		14'h311f:	ff_dbi <= 8'h00;
		14'h3120:	ff_dbi <= 8'h00;
		14'h3121:	ff_dbi <= 8'h00;
		14'h3122:	ff_dbi <= 8'h00;
		14'h3123:	ff_dbi <= 8'h00;
		14'h3124:	ff_dbi <= 8'h00;
		14'h3125:	ff_dbi <= 8'h00;
		14'h3126:	ff_dbi <= 8'h00;
		14'h3127:	ff_dbi <= 8'h00;
		14'h3128:	ff_dbi <= 8'h00;
		14'h3129:	ff_dbi <= 8'h00;
		14'h312a:	ff_dbi <= 8'h00;
		14'h312b:	ff_dbi <= 8'h00;
		14'h312c:	ff_dbi <= 8'h00;
		14'h312d:	ff_dbi <= 8'h00;
		14'h312e:	ff_dbi <= 8'h00;
		14'h312f:	ff_dbi <= 8'h00;
		14'h3130:	ff_dbi <= 8'h00;
		14'h3131:	ff_dbi <= 8'h00;
		14'h3132:	ff_dbi <= 8'h00;
		14'h3133:	ff_dbi <= 8'h00;
		14'h3134:	ff_dbi <= 8'h00;
		14'h3135:	ff_dbi <= 8'h00;
		14'h3136:	ff_dbi <= 8'h00;
		14'h3137:	ff_dbi <= 8'h00;
		14'h3138:	ff_dbi <= 8'h00;
		14'h3139:	ff_dbi <= 8'h00;
		14'h313a:	ff_dbi <= 8'h00;
		14'h313b:	ff_dbi <= 8'h00;
		14'h313c:	ff_dbi <= 8'h00;
		14'h313d:	ff_dbi <= 8'h00;
		14'h313e:	ff_dbi <= 8'h00;
		14'h313f:	ff_dbi <= 8'h00;
		14'h3140:	ff_dbi <= 8'h00;
		14'h3141:	ff_dbi <= 8'h00;
		14'h3142:	ff_dbi <= 8'h00;
		14'h3143:	ff_dbi <= 8'h00;
		14'h3144:	ff_dbi <= 8'h00;
		14'h3145:	ff_dbi <= 8'h00;
		14'h3146:	ff_dbi <= 8'h00;
		14'h3147:	ff_dbi <= 8'h00;
		14'h3148:	ff_dbi <= 8'h00;
		14'h3149:	ff_dbi <= 8'h00;
		14'h314a:	ff_dbi <= 8'h00;
		14'h314b:	ff_dbi <= 8'h00;
		14'h314c:	ff_dbi <= 8'h00;
		14'h314d:	ff_dbi <= 8'h00;
		14'h314e:	ff_dbi <= 8'h00;
		14'h314f:	ff_dbi <= 8'h00;
		14'h3150:	ff_dbi <= 8'h00;
		14'h3151:	ff_dbi <= 8'h00;
		14'h3152:	ff_dbi <= 8'h00;
		14'h3153:	ff_dbi <= 8'h00;
		14'h3154:	ff_dbi <= 8'h00;
		14'h3155:	ff_dbi <= 8'h00;
		14'h3156:	ff_dbi <= 8'h00;
		14'h3157:	ff_dbi <= 8'h00;
		14'h3158:	ff_dbi <= 8'h00;
		14'h3159:	ff_dbi <= 8'h00;
		14'h315a:	ff_dbi <= 8'h00;
		14'h315b:	ff_dbi <= 8'h00;
		14'h315c:	ff_dbi <= 8'h00;
		14'h315d:	ff_dbi <= 8'h00;
		14'h315e:	ff_dbi <= 8'h00;
		14'h315f:	ff_dbi <= 8'h00;
		14'h3160:	ff_dbi <= 8'h00;
		14'h3161:	ff_dbi <= 8'h00;
		14'h3162:	ff_dbi <= 8'h00;
		14'h3163:	ff_dbi <= 8'h00;
		14'h3164:	ff_dbi <= 8'h00;
		14'h3165:	ff_dbi <= 8'h00;
		14'h3166:	ff_dbi <= 8'h00;
		14'h3167:	ff_dbi <= 8'h00;
		14'h3168:	ff_dbi <= 8'h00;
		14'h3169:	ff_dbi <= 8'h00;
		14'h316a:	ff_dbi <= 8'h00;
		14'h316b:	ff_dbi <= 8'h00;
		14'h316c:	ff_dbi <= 8'h00;
		14'h316d:	ff_dbi <= 8'h00;
		14'h316e:	ff_dbi <= 8'h00;
		14'h316f:	ff_dbi <= 8'h00;
		14'h3170:	ff_dbi <= 8'h00;
		14'h3171:	ff_dbi <= 8'h00;
		14'h3172:	ff_dbi <= 8'h00;
		14'h3173:	ff_dbi <= 8'h00;
		14'h3174:	ff_dbi <= 8'h00;
		14'h3175:	ff_dbi <= 8'h00;
		14'h3176:	ff_dbi <= 8'h00;
		14'h3177:	ff_dbi <= 8'h00;
		14'h3178:	ff_dbi <= 8'h00;
		14'h3179:	ff_dbi <= 8'h00;
		14'h317a:	ff_dbi <= 8'h00;
		14'h317b:	ff_dbi <= 8'h00;
		14'h317c:	ff_dbi <= 8'h00;
		14'h317d:	ff_dbi <= 8'h00;
		14'h317e:	ff_dbi <= 8'h00;
		14'h317f:	ff_dbi <= 8'h00;
		14'h3180:	ff_dbi <= 8'h00;
		14'h3181:	ff_dbi <= 8'h00;
		14'h3182:	ff_dbi <= 8'h00;
		14'h3183:	ff_dbi <= 8'h00;
		14'h3184:	ff_dbi <= 8'h00;
		14'h3185:	ff_dbi <= 8'h00;
		14'h3186:	ff_dbi <= 8'h00;
		14'h3187:	ff_dbi <= 8'h00;
		14'h3188:	ff_dbi <= 8'h00;
		14'h3189:	ff_dbi <= 8'h00;
		14'h318a:	ff_dbi <= 8'h00;
		14'h318b:	ff_dbi <= 8'h00;
		14'h318c:	ff_dbi <= 8'h00;
		14'h318d:	ff_dbi <= 8'h00;
		14'h318e:	ff_dbi <= 8'h00;
		14'h318f:	ff_dbi <= 8'h00;
		14'h3190:	ff_dbi <= 8'h00;
		14'h3191:	ff_dbi <= 8'h00;
		14'h3192:	ff_dbi <= 8'h00;
		14'h3193:	ff_dbi <= 8'h00;
		14'h3194:	ff_dbi <= 8'h00;
		14'h3195:	ff_dbi <= 8'h00;
		14'h3196:	ff_dbi <= 8'h00;
		14'h3197:	ff_dbi <= 8'h00;
		14'h3198:	ff_dbi <= 8'h00;
		14'h3199:	ff_dbi <= 8'h00;
		14'h319a:	ff_dbi <= 8'h00;
		14'h319b:	ff_dbi <= 8'h00;
		14'h319c:	ff_dbi <= 8'h00;
		14'h319d:	ff_dbi <= 8'h00;
		14'h319e:	ff_dbi <= 8'h00;
		14'h319f:	ff_dbi <= 8'h00;
		14'h31a0:	ff_dbi <= 8'h00;
		14'h31a1:	ff_dbi <= 8'h00;
		14'h31a2:	ff_dbi <= 8'h00;
		14'h31a3:	ff_dbi <= 8'h00;
		14'h31a4:	ff_dbi <= 8'h00;
		14'h31a5:	ff_dbi <= 8'h00;
		14'h31a6:	ff_dbi <= 8'h00;
		14'h31a7:	ff_dbi <= 8'h00;
		14'h31a8:	ff_dbi <= 8'h00;
		14'h31a9:	ff_dbi <= 8'h00;
		14'h31aa:	ff_dbi <= 8'h00;
		14'h31ab:	ff_dbi <= 8'h00;
		14'h31ac:	ff_dbi <= 8'h00;
		14'h31ad:	ff_dbi <= 8'h00;
		14'h31ae:	ff_dbi <= 8'h00;
		14'h31af:	ff_dbi <= 8'h00;
		14'h31b0:	ff_dbi <= 8'h00;
		14'h31b1:	ff_dbi <= 8'h00;
		14'h31b2:	ff_dbi <= 8'h00;
		14'h31b3:	ff_dbi <= 8'h00;
		14'h31b4:	ff_dbi <= 8'h00;
		14'h31b5:	ff_dbi <= 8'h00;
		14'h31b6:	ff_dbi <= 8'h00;
		14'h31b7:	ff_dbi <= 8'h00;
		14'h31b8:	ff_dbi <= 8'h00;
		14'h31b9:	ff_dbi <= 8'h00;
		14'h31ba:	ff_dbi <= 8'h00;
		14'h31bb:	ff_dbi <= 8'h00;
		14'h31bc:	ff_dbi <= 8'h00;
		14'h31bd:	ff_dbi <= 8'h00;
		14'h31be:	ff_dbi <= 8'h00;
		14'h31bf:	ff_dbi <= 8'h00;
		14'h31c0:	ff_dbi <= 8'h00;
		14'h31c1:	ff_dbi <= 8'h00;
		14'h31c2:	ff_dbi <= 8'h00;
		14'h31c3:	ff_dbi <= 8'h00;
		14'h31c4:	ff_dbi <= 8'h00;
		14'h31c5:	ff_dbi <= 8'h00;
		14'h31c6:	ff_dbi <= 8'h00;
		14'h31c7:	ff_dbi <= 8'h00;
		14'h31c8:	ff_dbi <= 8'h00;
		14'h31c9:	ff_dbi <= 8'h00;
		14'h31ca:	ff_dbi <= 8'h00;
		14'h31cb:	ff_dbi <= 8'h00;
		14'h31cc:	ff_dbi <= 8'h00;
		14'h31cd:	ff_dbi <= 8'h00;
		14'h31ce:	ff_dbi <= 8'h00;
		14'h31cf:	ff_dbi <= 8'h00;
		14'h31d0:	ff_dbi <= 8'h00;
		14'h31d1:	ff_dbi <= 8'h00;
		14'h31d2:	ff_dbi <= 8'h00;
		14'h31d3:	ff_dbi <= 8'h00;
		14'h31d4:	ff_dbi <= 8'h00;
		14'h31d5:	ff_dbi <= 8'h00;
		14'h31d6:	ff_dbi <= 8'h00;
		14'h31d7:	ff_dbi <= 8'h00;
		14'h31d8:	ff_dbi <= 8'h00;
		14'h31d9:	ff_dbi <= 8'h00;
		14'h31da:	ff_dbi <= 8'h00;
		14'h31db:	ff_dbi <= 8'h00;
		14'h31dc:	ff_dbi <= 8'h00;
		14'h31dd:	ff_dbi <= 8'h00;
		14'h31de:	ff_dbi <= 8'h00;
		14'h31df:	ff_dbi <= 8'h00;
		14'h31e0:	ff_dbi <= 8'h00;
		14'h31e1:	ff_dbi <= 8'h00;
		14'h31e2:	ff_dbi <= 8'h00;
		14'h31e3:	ff_dbi <= 8'h00;
		14'h31e4:	ff_dbi <= 8'h00;
		14'h31e5:	ff_dbi <= 8'h00;
		14'h31e6:	ff_dbi <= 8'h00;
		14'h31e7:	ff_dbi <= 8'h00;
		14'h31e8:	ff_dbi <= 8'h00;
		14'h31e9:	ff_dbi <= 8'h00;
		14'h31ea:	ff_dbi <= 8'h00;
		14'h31eb:	ff_dbi <= 8'h00;
		14'h31ec:	ff_dbi <= 8'h00;
		14'h31ed:	ff_dbi <= 8'h00;
		14'h31ee:	ff_dbi <= 8'h00;
		14'h31ef:	ff_dbi <= 8'h00;
		14'h31f0:	ff_dbi <= 8'h00;
		14'h31f1:	ff_dbi <= 8'h00;
		14'h31f2:	ff_dbi <= 8'h00;
		14'h31f3:	ff_dbi <= 8'h00;
		14'h31f4:	ff_dbi <= 8'h00;
		14'h31f5:	ff_dbi <= 8'h00;
		14'h31f6:	ff_dbi <= 8'h00;
		14'h31f7:	ff_dbi <= 8'h00;
		14'h31f8:	ff_dbi <= 8'h00;
		14'h31f9:	ff_dbi <= 8'h00;
		14'h31fa:	ff_dbi <= 8'h00;
		14'h31fb:	ff_dbi <= 8'h00;
		14'h31fc:	ff_dbi <= 8'h00;
		14'h31fd:	ff_dbi <= 8'h00;
		14'h31fe:	ff_dbi <= 8'h00;
		14'h31ff:	ff_dbi <= 8'h00;
		14'h3200:	ff_dbi <= 8'h00;
		14'h3201:	ff_dbi <= 8'h00;
		14'h3202:	ff_dbi <= 8'h00;
		14'h3203:	ff_dbi <= 8'h00;
		14'h3204:	ff_dbi <= 8'h00;
		14'h3205:	ff_dbi <= 8'h00;
		14'h3206:	ff_dbi <= 8'h00;
		14'h3207:	ff_dbi <= 8'h00;
		14'h3208:	ff_dbi <= 8'h00;
		14'h3209:	ff_dbi <= 8'h00;
		14'h320a:	ff_dbi <= 8'h00;
		14'h320b:	ff_dbi <= 8'h00;
		14'h320c:	ff_dbi <= 8'h00;
		14'h320d:	ff_dbi <= 8'h00;
		14'h320e:	ff_dbi <= 8'h00;
		14'h320f:	ff_dbi <= 8'h00;
		14'h3210:	ff_dbi <= 8'h00;
		14'h3211:	ff_dbi <= 8'h00;
		14'h3212:	ff_dbi <= 8'h00;
		14'h3213:	ff_dbi <= 8'h00;
		14'h3214:	ff_dbi <= 8'h00;
		14'h3215:	ff_dbi <= 8'h00;
		14'h3216:	ff_dbi <= 8'h00;
		14'h3217:	ff_dbi <= 8'h00;
		14'h3218:	ff_dbi <= 8'h00;
		14'h3219:	ff_dbi <= 8'h00;
		14'h321a:	ff_dbi <= 8'h00;
		14'h321b:	ff_dbi <= 8'h00;
		14'h321c:	ff_dbi <= 8'h00;
		14'h321d:	ff_dbi <= 8'h00;
		14'h321e:	ff_dbi <= 8'h00;
		14'h321f:	ff_dbi <= 8'h00;
		14'h3220:	ff_dbi <= 8'h00;
		14'h3221:	ff_dbi <= 8'h00;
		14'h3222:	ff_dbi <= 8'h00;
		14'h3223:	ff_dbi <= 8'h00;
		14'h3224:	ff_dbi <= 8'h00;
		14'h3225:	ff_dbi <= 8'h00;
		14'h3226:	ff_dbi <= 8'h00;
		14'h3227:	ff_dbi <= 8'h00;
		14'h3228:	ff_dbi <= 8'h00;
		14'h3229:	ff_dbi <= 8'h00;
		14'h322a:	ff_dbi <= 8'h00;
		14'h322b:	ff_dbi <= 8'h00;
		14'h322c:	ff_dbi <= 8'h00;
		14'h322d:	ff_dbi <= 8'h00;
		14'h322e:	ff_dbi <= 8'h00;
		14'h322f:	ff_dbi <= 8'h00;
		14'h3230:	ff_dbi <= 8'h00;
		14'h3231:	ff_dbi <= 8'h00;
		14'h3232:	ff_dbi <= 8'h00;
		14'h3233:	ff_dbi <= 8'h00;
		14'h3234:	ff_dbi <= 8'h00;
		14'h3235:	ff_dbi <= 8'h00;
		14'h3236:	ff_dbi <= 8'h00;
		14'h3237:	ff_dbi <= 8'h00;
		14'h3238:	ff_dbi <= 8'h00;
		14'h3239:	ff_dbi <= 8'h00;
		14'h323a:	ff_dbi <= 8'h00;
		14'h323b:	ff_dbi <= 8'h00;
		14'h323c:	ff_dbi <= 8'h00;
		14'h323d:	ff_dbi <= 8'h00;
		14'h323e:	ff_dbi <= 8'h00;
		14'h323f:	ff_dbi <= 8'h00;
		14'h3240:	ff_dbi <= 8'h00;
		14'h3241:	ff_dbi <= 8'h00;
		14'h3242:	ff_dbi <= 8'h00;
		14'h3243:	ff_dbi <= 8'h00;
		14'h3244:	ff_dbi <= 8'h00;
		14'h3245:	ff_dbi <= 8'h00;
		14'h3246:	ff_dbi <= 8'h00;
		14'h3247:	ff_dbi <= 8'h00;
		14'h3248:	ff_dbi <= 8'h00;
		14'h3249:	ff_dbi <= 8'h00;
		14'h324a:	ff_dbi <= 8'h00;
		14'h324b:	ff_dbi <= 8'h00;
		14'h324c:	ff_dbi <= 8'h00;
		14'h324d:	ff_dbi <= 8'h00;
		14'h324e:	ff_dbi <= 8'h00;
		14'h324f:	ff_dbi <= 8'h00;
		14'h3250:	ff_dbi <= 8'h00;
		14'h3251:	ff_dbi <= 8'h00;
		14'h3252:	ff_dbi <= 8'h00;
		14'h3253:	ff_dbi <= 8'h00;
		14'h3254:	ff_dbi <= 8'h00;
		14'h3255:	ff_dbi <= 8'h00;
		14'h3256:	ff_dbi <= 8'h00;
		14'h3257:	ff_dbi <= 8'h00;
		14'h3258:	ff_dbi <= 8'h00;
		14'h3259:	ff_dbi <= 8'h00;
		14'h325a:	ff_dbi <= 8'h00;
		14'h325b:	ff_dbi <= 8'h00;
		14'h325c:	ff_dbi <= 8'h00;
		14'h325d:	ff_dbi <= 8'h00;
		14'h325e:	ff_dbi <= 8'h00;
		14'h325f:	ff_dbi <= 8'h00;
		14'h3260:	ff_dbi <= 8'h00;
		14'h3261:	ff_dbi <= 8'h00;
		14'h3262:	ff_dbi <= 8'h00;
		14'h3263:	ff_dbi <= 8'h00;
		14'h3264:	ff_dbi <= 8'h00;
		14'h3265:	ff_dbi <= 8'h00;
		14'h3266:	ff_dbi <= 8'h00;
		14'h3267:	ff_dbi <= 8'h00;
		14'h3268:	ff_dbi <= 8'h00;
		14'h3269:	ff_dbi <= 8'h00;
		14'h326a:	ff_dbi <= 8'h00;
		14'h326b:	ff_dbi <= 8'h00;
		14'h326c:	ff_dbi <= 8'h00;
		14'h326d:	ff_dbi <= 8'h00;
		14'h326e:	ff_dbi <= 8'h00;
		14'h326f:	ff_dbi <= 8'h00;
		14'h3270:	ff_dbi <= 8'h00;
		14'h3271:	ff_dbi <= 8'h00;
		14'h3272:	ff_dbi <= 8'h00;
		14'h3273:	ff_dbi <= 8'h00;
		14'h3274:	ff_dbi <= 8'h00;
		14'h3275:	ff_dbi <= 8'h00;
		14'h3276:	ff_dbi <= 8'h00;
		14'h3277:	ff_dbi <= 8'h00;
		14'h3278:	ff_dbi <= 8'h00;
		14'h3279:	ff_dbi <= 8'h00;
		14'h327a:	ff_dbi <= 8'h00;
		14'h327b:	ff_dbi <= 8'h00;
		14'h327c:	ff_dbi <= 8'h00;
		14'h327d:	ff_dbi <= 8'h00;
		14'h327e:	ff_dbi <= 8'h00;
		14'h327f:	ff_dbi <= 8'h00;
		14'h3280:	ff_dbi <= 8'h00;
		14'h3281:	ff_dbi <= 8'h00;
		14'h3282:	ff_dbi <= 8'h00;
		14'h3283:	ff_dbi <= 8'h00;
		14'h3284:	ff_dbi <= 8'h00;
		14'h3285:	ff_dbi <= 8'h00;
		14'h3286:	ff_dbi <= 8'h00;
		14'h3287:	ff_dbi <= 8'h00;
		14'h3288:	ff_dbi <= 8'h00;
		14'h3289:	ff_dbi <= 8'h00;
		14'h328a:	ff_dbi <= 8'h00;
		14'h328b:	ff_dbi <= 8'h00;
		14'h328c:	ff_dbi <= 8'h00;
		14'h328d:	ff_dbi <= 8'h00;
		14'h328e:	ff_dbi <= 8'h00;
		14'h328f:	ff_dbi <= 8'h00;
		14'h3290:	ff_dbi <= 8'h00;
		14'h3291:	ff_dbi <= 8'h00;
		14'h3292:	ff_dbi <= 8'h00;
		14'h3293:	ff_dbi <= 8'h00;
		14'h3294:	ff_dbi <= 8'h00;
		14'h3295:	ff_dbi <= 8'h00;
		14'h3296:	ff_dbi <= 8'h00;
		14'h3297:	ff_dbi <= 8'h00;
		14'h3298:	ff_dbi <= 8'h00;
		14'h3299:	ff_dbi <= 8'h00;
		14'h329a:	ff_dbi <= 8'h00;
		14'h329b:	ff_dbi <= 8'h00;
		14'h329c:	ff_dbi <= 8'h00;
		14'h329d:	ff_dbi <= 8'h00;
		14'h329e:	ff_dbi <= 8'h00;
		14'h329f:	ff_dbi <= 8'h00;
		14'h32a0:	ff_dbi <= 8'h00;
		14'h32a1:	ff_dbi <= 8'h00;
		14'h32a2:	ff_dbi <= 8'h00;
		14'h32a3:	ff_dbi <= 8'h00;
		14'h32a4:	ff_dbi <= 8'h00;
		14'h32a5:	ff_dbi <= 8'h00;
		14'h32a6:	ff_dbi <= 8'h00;
		14'h32a7:	ff_dbi <= 8'h00;
		14'h32a8:	ff_dbi <= 8'h00;
		14'h32a9:	ff_dbi <= 8'h00;
		14'h32aa:	ff_dbi <= 8'h00;
		14'h32ab:	ff_dbi <= 8'h00;
		14'h32ac:	ff_dbi <= 8'h00;
		14'h32ad:	ff_dbi <= 8'h00;
		14'h32ae:	ff_dbi <= 8'h00;
		14'h32af:	ff_dbi <= 8'h00;
		14'h32b0:	ff_dbi <= 8'h00;
		14'h32b1:	ff_dbi <= 8'h00;
		14'h32b2:	ff_dbi <= 8'h00;
		14'h32b3:	ff_dbi <= 8'h00;
		14'h32b4:	ff_dbi <= 8'h00;
		14'h32b5:	ff_dbi <= 8'h00;
		14'h32b6:	ff_dbi <= 8'h00;
		14'h32b7:	ff_dbi <= 8'h00;
		14'h32b8:	ff_dbi <= 8'h00;
		14'h32b9:	ff_dbi <= 8'h00;
		14'h32ba:	ff_dbi <= 8'h00;
		14'h32bb:	ff_dbi <= 8'h00;
		14'h32bc:	ff_dbi <= 8'h00;
		14'h32bd:	ff_dbi <= 8'h00;
		14'h32be:	ff_dbi <= 8'h00;
		14'h32bf:	ff_dbi <= 8'h00;
		14'h32c0:	ff_dbi <= 8'h00;
		14'h32c1:	ff_dbi <= 8'h00;
		14'h32c2:	ff_dbi <= 8'h00;
		14'h32c3:	ff_dbi <= 8'h00;
		14'h32c4:	ff_dbi <= 8'h00;
		14'h32c5:	ff_dbi <= 8'h00;
		14'h32c6:	ff_dbi <= 8'h00;
		14'h32c7:	ff_dbi <= 8'h00;
		14'h32c8:	ff_dbi <= 8'h00;
		14'h32c9:	ff_dbi <= 8'h00;
		14'h32ca:	ff_dbi <= 8'h00;
		14'h32cb:	ff_dbi <= 8'h00;
		14'h32cc:	ff_dbi <= 8'h00;
		14'h32cd:	ff_dbi <= 8'h00;
		14'h32ce:	ff_dbi <= 8'h00;
		14'h32cf:	ff_dbi <= 8'h00;
		14'h32d0:	ff_dbi <= 8'h00;
		14'h32d1:	ff_dbi <= 8'h00;
		14'h32d2:	ff_dbi <= 8'h00;
		14'h32d3:	ff_dbi <= 8'h00;
		14'h32d4:	ff_dbi <= 8'h00;
		14'h32d5:	ff_dbi <= 8'h00;
		14'h32d6:	ff_dbi <= 8'h00;
		14'h32d7:	ff_dbi <= 8'h00;
		14'h32d8:	ff_dbi <= 8'h00;
		14'h32d9:	ff_dbi <= 8'h00;
		14'h32da:	ff_dbi <= 8'h00;
		14'h32db:	ff_dbi <= 8'h00;
		14'h32dc:	ff_dbi <= 8'h00;
		14'h32dd:	ff_dbi <= 8'h00;
		14'h32de:	ff_dbi <= 8'h00;
		14'h32df:	ff_dbi <= 8'h00;
		14'h32e0:	ff_dbi <= 8'h00;
		14'h32e1:	ff_dbi <= 8'h00;
		14'h32e2:	ff_dbi <= 8'h00;
		14'h32e3:	ff_dbi <= 8'h00;
		14'h32e4:	ff_dbi <= 8'h00;
		14'h32e5:	ff_dbi <= 8'h00;
		14'h32e6:	ff_dbi <= 8'h00;
		14'h32e7:	ff_dbi <= 8'h00;
		14'h32e8:	ff_dbi <= 8'h00;
		14'h32e9:	ff_dbi <= 8'h00;
		14'h32ea:	ff_dbi <= 8'h00;
		14'h32eb:	ff_dbi <= 8'h00;
		14'h32ec:	ff_dbi <= 8'h00;
		14'h32ed:	ff_dbi <= 8'h00;
		14'h32ee:	ff_dbi <= 8'h00;
		14'h32ef:	ff_dbi <= 8'h00;
		14'h32f0:	ff_dbi <= 8'h00;
		14'h32f1:	ff_dbi <= 8'h00;
		14'h32f2:	ff_dbi <= 8'h00;
		14'h32f3:	ff_dbi <= 8'h00;
		14'h32f4:	ff_dbi <= 8'h00;
		14'h32f5:	ff_dbi <= 8'h00;
		14'h32f6:	ff_dbi <= 8'h00;
		14'h32f7:	ff_dbi <= 8'h00;
		14'h32f8:	ff_dbi <= 8'h00;
		14'h32f9:	ff_dbi <= 8'h00;
		14'h32fa:	ff_dbi <= 8'h00;
		14'h32fb:	ff_dbi <= 8'h00;
		14'h32fc:	ff_dbi <= 8'h00;
		14'h32fd:	ff_dbi <= 8'h00;
		14'h32fe:	ff_dbi <= 8'h00;
		14'h32ff:	ff_dbi <= 8'h00;
		14'h3300:	ff_dbi <= 8'h00;
		14'h3301:	ff_dbi <= 8'h00;
		14'h3302:	ff_dbi <= 8'h00;
		14'h3303:	ff_dbi <= 8'h00;
		14'h3304:	ff_dbi <= 8'h00;
		14'h3305:	ff_dbi <= 8'h00;
		14'h3306:	ff_dbi <= 8'h00;
		14'h3307:	ff_dbi <= 8'h00;
		14'h3308:	ff_dbi <= 8'h00;
		14'h3309:	ff_dbi <= 8'h00;
		14'h330a:	ff_dbi <= 8'h00;
		14'h330b:	ff_dbi <= 8'h00;
		14'h330c:	ff_dbi <= 8'h00;
		14'h330d:	ff_dbi <= 8'h00;
		14'h330e:	ff_dbi <= 8'h00;
		14'h330f:	ff_dbi <= 8'h00;
		14'h3310:	ff_dbi <= 8'h00;
		14'h3311:	ff_dbi <= 8'h00;
		14'h3312:	ff_dbi <= 8'h00;
		14'h3313:	ff_dbi <= 8'h00;
		14'h3314:	ff_dbi <= 8'h00;
		14'h3315:	ff_dbi <= 8'h00;
		14'h3316:	ff_dbi <= 8'h00;
		14'h3317:	ff_dbi <= 8'h00;
		14'h3318:	ff_dbi <= 8'h00;
		14'h3319:	ff_dbi <= 8'h00;
		14'h331a:	ff_dbi <= 8'h00;
		14'h331b:	ff_dbi <= 8'h00;
		14'h331c:	ff_dbi <= 8'h00;
		14'h331d:	ff_dbi <= 8'h00;
		14'h331e:	ff_dbi <= 8'h00;
		14'h331f:	ff_dbi <= 8'h00;
		14'h3320:	ff_dbi <= 8'h00;
		14'h3321:	ff_dbi <= 8'h00;
		14'h3322:	ff_dbi <= 8'h00;
		14'h3323:	ff_dbi <= 8'h00;
		14'h3324:	ff_dbi <= 8'h00;
		14'h3325:	ff_dbi <= 8'h00;
		14'h3326:	ff_dbi <= 8'h00;
		14'h3327:	ff_dbi <= 8'h00;
		14'h3328:	ff_dbi <= 8'h00;
		14'h3329:	ff_dbi <= 8'h00;
		14'h332a:	ff_dbi <= 8'h00;
		14'h332b:	ff_dbi <= 8'h00;
		14'h332c:	ff_dbi <= 8'h00;
		14'h332d:	ff_dbi <= 8'h00;
		14'h332e:	ff_dbi <= 8'h00;
		14'h332f:	ff_dbi <= 8'h00;
		14'h3330:	ff_dbi <= 8'h00;
		14'h3331:	ff_dbi <= 8'h00;
		14'h3332:	ff_dbi <= 8'h00;
		14'h3333:	ff_dbi <= 8'h00;
		14'h3334:	ff_dbi <= 8'h00;
		14'h3335:	ff_dbi <= 8'h00;
		14'h3336:	ff_dbi <= 8'h00;
		14'h3337:	ff_dbi <= 8'h00;
		14'h3338:	ff_dbi <= 8'h00;
		14'h3339:	ff_dbi <= 8'h00;
		14'h333a:	ff_dbi <= 8'h00;
		14'h333b:	ff_dbi <= 8'h00;
		14'h333c:	ff_dbi <= 8'h00;
		14'h333d:	ff_dbi <= 8'h00;
		14'h333e:	ff_dbi <= 8'h00;
		14'h333f:	ff_dbi <= 8'h00;
		14'h3340:	ff_dbi <= 8'h00;
		14'h3341:	ff_dbi <= 8'h00;
		14'h3342:	ff_dbi <= 8'h00;
		14'h3343:	ff_dbi <= 8'h00;
		14'h3344:	ff_dbi <= 8'h00;
		14'h3345:	ff_dbi <= 8'h00;
		14'h3346:	ff_dbi <= 8'h00;
		14'h3347:	ff_dbi <= 8'h00;
		14'h3348:	ff_dbi <= 8'h00;
		14'h3349:	ff_dbi <= 8'h00;
		14'h334a:	ff_dbi <= 8'h00;
		14'h334b:	ff_dbi <= 8'h00;
		14'h334c:	ff_dbi <= 8'h00;
		14'h334d:	ff_dbi <= 8'h00;
		14'h334e:	ff_dbi <= 8'h00;
		14'h334f:	ff_dbi <= 8'h00;
		14'h3350:	ff_dbi <= 8'h00;
		14'h3351:	ff_dbi <= 8'h00;
		14'h3352:	ff_dbi <= 8'h00;
		14'h3353:	ff_dbi <= 8'h00;
		14'h3354:	ff_dbi <= 8'h00;
		14'h3355:	ff_dbi <= 8'h00;
		14'h3356:	ff_dbi <= 8'h00;
		14'h3357:	ff_dbi <= 8'h00;
		14'h3358:	ff_dbi <= 8'h00;
		14'h3359:	ff_dbi <= 8'h00;
		14'h335a:	ff_dbi <= 8'h00;
		14'h335b:	ff_dbi <= 8'h00;
		14'h335c:	ff_dbi <= 8'h00;
		14'h335d:	ff_dbi <= 8'h00;
		14'h335e:	ff_dbi <= 8'h00;
		14'h335f:	ff_dbi <= 8'h00;
		14'h3360:	ff_dbi <= 8'h00;
		14'h3361:	ff_dbi <= 8'h00;
		14'h3362:	ff_dbi <= 8'h00;
		14'h3363:	ff_dbi <= 8'h00;
		14'h3364:	ff_dbi <= 8'h00;
		14'h3365:	ff_dbi <= 8'h00;
		14'h3366:	ff_dbi <= 8'h00;
		14'h3367:	ff_dbi <= 8'h00;
		14'h3368:	ff_dbi <= 8'h00;
		14'h3369:	ff_dbi <= 8'h00;
		14'h336a:	ff_dbi <= 8'h00;
		14'h336b:	ff_dbi <= 8'h00;
		14'h336c:	ff_dbi <= 8'h00;
		14'h336d:	ff_dbi <= 8'h00;
		14'h336e:	ff_dbi <= 8'h00;
		14'h336f:	ff_dbi <= 8'h00;
		14'h3370:	ff_dbi <= 8'h00;
		14'h3371:	ff_dbi <= 8'h00;
		14'h3372:	ff_dbi <= 8'h00;
		14'h3373:	ff_dbi <= 8'h00;
		14'h3374:	ff_dbi <= 8'h00;
		14'h3375:	ff_dbi <= 8'h00;
		14'h3376:	ff_dbi <= 8'h00;
		14'h3377:	ff_dbi <= 8'h00;
		14'h3378:	ff_dbi <= 8'h00;
		14'h3379:	ff_dbi <= 8'h00;
		14'h337a:	ff_dbi <= 8'h00;
		14'h337b:	ff_dbi <= 8'h00;
		14'h337c:	ff_dbi <= 8'h00;
		14'h337d:	ff_dbi <= 8'h00;
		14'h337e:	ff_dbi <= 8'h00;
		14'h337f:	ff_dbi <= 8'h00;
		14'h3380:	ff_dbi <= 8'h00;
		14'h3381:	ff_dbi <= 8'h00;
		14'h3382:	ff_dbi <= 8'h00;
		14'h3383:	ff_dbi <= 8'h00;
		14'h3384:	ff_dbi <= 8'h00;
		14'h3385:	ff_dbi <= 8'h00;
		14'h3386:	ff_dbi <= 8'h00;
		14'h3387:	ff_dbi <= 8'h00;
		14'h3388:	ff_dbi <= 8'h00;
		14'h3389:	ff_dbi <= 8'h00;
		14'h338a:	ff_dbi <= 8'h00;
		14'h338b:	ff_dbi <= 8'h00;
		14'h338c:	ff_dbi <= 8'h00;
		14'h338d:	ff_dbi <= 8'h00;
		14'h338e:	ff_dbi <= 8'h00;
		14'h338f:	ff_dbi <= 8'h00;
		14'h3390:	ff_dbi <= 8'h00;
		14'h3391:	ff_dbi <= 8'h00;
		14'h3392:	ff_dbi <= 8'h00;
		14'h3393:	ff_dbi <= 8'h00;
		14'h3394:	ff_dbi <= 8'h00;
		14'h3395:	ff_dbi <= 8'h00;
		14'h3396:	ff_dbi <= 8'h00;
		14'h3397:	ff_dbi <= 8'h00;
		14'h3398:	ff_dbi <= 8'h00;
		14'h3399:	ff_dbi <= 8'h00;
		14'h339a:	ff_dbi <= 8'h00;
		14'h339b:	ff_dbi <= 8'h00;
		14'h339c:	ff_dbi <= 8'h00;
		14'h339d:	ff_dbi <= 8'h00;
		14'h339e:	ff_dbi <= 8'h00;
		14'h339f:	ff_dbi <= 8'h00;
		14'h33a0:	ff_dbi <= 8'h00;
		14'h33a1:	ff_dbi <= 8'h00;
		14'h33a2:	ff_dbi <= 8'h00;
		14'h33a3:	ff_dbi <= 8'h00;
		14'h33a4:	ff_dbi <= 8'h00;
		14'h33a5:	ff_dbi <= 8'h00;
		14'h33a6:	ff_dbi <= 8'h00;
		14'h33a7:	ff_dbi <= 8'h00;
		14'h33a8:	ff_dbi <= 8'h00;
		14'h33a9:	ff_dbi <= 8'h00;
		14'h33aa:	ff_dbi <= 8'h00;
		14'h33ab:	ff_dbi <= 8'h00;
		14'h33ac:	ff_dbi <= 8'h00;
		14'h33ad:	ff_dbi <= 8'h00;
		14'h33ae:	ff_dbi <= 8'h00;
		14'h33af:	ff_dbi <= 8'h00;
		14'h33b0:	ff_dbi <= 8'h00;
		14'h33b1:	ff_dbi <= 8'h00;
		14'h33b2:	ff_dbi <= 8'h00;
		14'h33b3:	ff_dbi <= 8'h00;
		14'h33b4:	ff_dbi <= 8'h00;
		14'h33b5:	ff_dbi <= 8'h00;
		14'h33b6:	ff_dbi <= 8'h00;
		14'h33b7:	ff_dbi <= 8'h00;
		14'h33b8:	ff_dbi <= 8'h00;
		14'h33b9:	ff_dbi <= 8'h00;
		14'h33ba:	ff_dbi <= 8'h00;
		14'h33bb:	ff_dbi <= 8'h00;
		14'h33bc:	ff_dbi <= 8'h00;
		14'h33bd:	ff_dbi <= 8'h00;
		14'h33be:	ff_dbi <= 8'h00;
		14'h33bf:	ff_dbi <= 8'h00;
		14'h33c0:	ff_dbi <= 8'h00;
		14'h33c1:	ff_dbi <= 8'h00;
		14'h33c2:	ff_dbi <= 8'h00;
		14'h33c3:	ff_dbi <= 8'h00;
		14'h33c4:	ff_dbi <= 8'h00;
		14'h33c5:	ff_dbi <= 8'h00;
		14'h33c6:	ff_dbi <= 8'h00;
		14'h33c7:	ff_dbi <= 8'h00;
		14'h33c8:	ff_dbi <= 8'h00;
		14'h33c9:	ff_dbi <= 8'h00;
		14'h33ca:	ff_dbi <= 8'h00;
		14'h33cb:	ff_dbi <= 8'h00;
		14'h33cc:	ff_dbi <= 8'h00;
		14'h33cd:	ff_dbi <= 8'h00;
		14'h33ce:	ff_dbi <= 8'h00;
		14'h33cf:	ff_dbi <= 8'h00;
		14'h33d0:	ff_dbi <= 8'h00;
		14'h33d1:	ff_dbi <= 8'h00;
		14'h33d2:	ff_dbi <= 8'h00;
		14'h33d3:	ff_dbi <= 8'h00;
		14'h33d4:	ff_dbi <= 8'h00;
		14'h33d5:	ff_dbi <= 8'h00;
		14'h33d6:	ff_dbi <= 8'h00;
		14'h33d7:	ff_dbi <= 8'h00;
		14'h33d8:	ff_dbi <= 8'h00;
		14'h33d9:	ff_dbi <= 8'h00;
		14'h33da:	ff_dbi <= 8'h00;
		14'h33db:	ff_dbi <= 8'h00;
		14'h33dc:	ff_dbi <= 8'h00;
		14'h33dd:	ff_dbi <= 8'h00;
		14'h33de:	ff_dbi <= 8'h00;
		14'h33df:	ff_dbi <= 8'h00;
		14'h33e0:	ff_dbi <= 8'h00;
		14'h33e1:	ff_dbi <= 8'h00;
		14'h33e2:	ff_dbi <= 8'h00;
		14'h33e3:	ff_dbi <= 8'h00;
		14'h33e4:	ff_dbi <= 8'h00;
		14'h33e5:	ff_dbi <= 8'h00;
		14'h33e6:	ff_dbi <= 8'h00;
		14'h33e7:	ff_dbi <= 8'h00;
		14'h33e8:	ff_dbi <= 8'h00;
		14'h33e9:	ff_dbi <= 8'h00;
		14'h33ea:	ff_dbi <= 8'h00;
		14'h33eb:	ff_dbi <= 8'h00;
		14'h33ec:	ff_dbi <= 8'h00;
		14'h33ed:	ff_dbi <= 8'h00;
		14'h33ee:	ff_dbi <= 8'h00;
		14'h33ef:	ff_dbi <= 8'h00;
		14'h33f0:	ff_dbi <= 8'h00;
		14'h33f1:	ff_dbi <= 8'h00;
		14'h33f2:	ff_dbi <= 8'h00;
		14'h33f3:	ff_dbi <= 8'h00;
		14'h33f4:	ff_dbi <= 8'h00;
		14'h33f5:	ff_dbi <= 8'h00;
		14'h33f6:	ff_dbi <= 8'h00;
		14'h33f7:	ff_dbi <= 8'h00;
		14'h33f8:	ff_dbi <= 8'h00;
		14'h33f9:	ff_dbi <= 8'h00;
		14'h33fa:	ff_dbi <= 8'h00;
		14'h33fb:	ff_dbi <= 8'h00;
		14'h33fc:	ff_dbi <= 8'h00;
		14'h33fd:	ff_dbi <= 8'h00;
		14'h33fe:	ff_dbi <= 8'h00;
		14'h33ff:	ff_dbi <= 8'h00;
		14'h3400:	ff_dbi <= 8'h00;
		14'h3401:	ff_dbi <= 8'h00;
		14'h3402:	ff_dbi <= 8'h00;
		14'h3403:	ff_dbi <= 8'h00;
		14'h3404:	ff_dbi <= 8'h00;
		14'h3405:	ff_dbi <= 8'h00;
		14'h3406:	ff_dbi <= 8'h00;
		14'h3407:	ff_dbi <= 8'h00;
		14'h3408:	ff_dbi <= 8'h00;
		14'h3409:	ff_dbi <= 8'h00;
		14'h340a:	ff_dbi <= 8'h00;
		14'h340b:	ff_dbi <= 8'h00;
		14'h340c:	ff_dbi <= 8'h00;
		14'h340d:	ff_dbi <= 8'h00;
		14'h340e:	ff_dbi <= 8'h00;
		14'h340f:	ff_dbi <= 8'h00;
		14'h3410:	ff_dbi <= 8'h00;
		14'h3411:	ff_dbi <= 8'h00;
		14'h3412:	ff_dbi <= 8'h00;
		14'h3413:	ff_dbi <= 8'h00;
		14'h3414:	ff_dbi <= 8'h00;
		14'h3415:	ff_dbi <= 8'h00;
		14'h3416:	ff_dbi <= 8'h00;
		14'h3417:	ff_dbi <= 8'h00;
		14'h3418:	ff_dbi <= 8'h00;
		14'h3419:	ff_dbi <= 8'h00;
		14'h341a:	ff_dbi <= 8'h00;
		14'h341b:	ff_dbi <= 8'h00;
		14'h341c:	ff_dbi <= 8'h00;
		14'h341d:	ff_dbi <= 8'h00;
		14'h341e:	ff_dbi <= 8'h00;
		14'h341f:	ff_dbi <= 8'h00;
		14'h3420:	ff_dbi <= 8'h00;
		14'h3421:	ff_dbi <= 8'h00;
		14'h3422:	ff_dbi <= 8'h00;
		14'h3423:	ff_dbi <= 8'h00;
		14'h3424:	ff_dbi <= 8'h00;
		14'h3425:	ff_dbi <= 8'h00;
		14'h3426:	ff_dbi <= 8'h00;
		14'h3427:	ff_dbi <= 8'h00;
		14'h3428:	ff_dbi <= 8'h00;
		14'h3429:	ff_dbi <= 8'h00;
		14'h342a:	ff_dbi <= 8'h00;
		14'h342b:	ff_dbi <= 8'h00;
		14'h342c:	ff_dbi <= 8'h00;
		14'h342d:	ff_dbi <= 8'h00;
		14'h342e:	ff_dbi <= 8'h00;
		14'h342f:	ff_dbi <= 8'h00;
		14'h3430:	ff_dbi <= 8'h00;
		14'h3431:	ff_dbi <= 8'h00;
		14'h3432:	ff_dbi <= 8'h00;
		14'h3433:	ff_dbi <= 8'h00;
		14'h3434:	ff_dbi <= 8'h00;
		14'h3435:	ff_dbi <= 8'h00;
		14'h3436:	ff_dbi <= 8'h00;
		14'h3437:	ff_dbi <= 8'h00;
		14'h3438:	ff_dbi <= 8'h00;
		14'h3439:	ff_dbi <= 8'h00;
		14'h343a:	ff_dbi <= 8'h00;
		14'h343b:	ff_dbi <= 8'h00;
		14'h343c:	ff_dbi <= 8'h00;
		14'h343d:	ff_dbi <= 8'h00;
		14'h343e:	ff_dbi <= 8'h00;
		14'h343f:	ff_dbi <= 8'h00;
		14'h3440:	ff_dbi <= 8'h00;
		14'h3441:	ff_dbi <= 8'h00;
		14'h3442:	ff_dbi <= 8'h00;
		14'h3443:	ff_dbi <= 8'h00;
		14'h3444:	ff_dbi <= 8'h00;
		14'h3445:	ff_dbi <= 8'h00;
		14'h3446:	ff_dbi <= 8'h00;
		14'h3447:	ff_dbi <= 8'h00;
		14'h3448:	ff_dbi <= 8'h00;
		14'h3449:	ff_dbi <= 8'h00;
		14'h344a:	ff_dbi <= 8'h00;
		14'h344b:	ff_dbi <= 8'h00;
		14'h344c:	ff_dbi <= 8'h00;
		14'h344d:	ff_dbi <= 8'h00;
		14'h344e:	ff_dbi <= 8'h00;
		14'h344f:	ff_dbi <= 8'h00;
		14'h3450:	ff_dbi <= 8'h00;
		14'h3451:	ff_dbi <= 8'h00;
		14'h3452:	ff_dbi <= 8'h00;
		14'h3453:	ff_dbi <= 8'h00;
		14'h3454:	ff_dbi <= 8'h00;
		14'h3455:	ff_dbi <= 8'h00;
		14'h3456:	ff_dbi <= 8'h00;
		14'h3457:	ff_dbi <= 8'h00;
		14'h3458:	ff_dbi <= 8'h00;
		14'h3459:	ff_dbi <= 8'h00;
		14'h345a:	ff_dbi <= 8'h00;
		14'h345b:	ff_dbi <= 8'h00;
		14'h345c:	ff_dbi <= 8'h00;
		14'h345d:	ff_dbi <= 8'h00;
		14'h345e:	ff_dbi <= 8'h00;
		14'h345f:	ff_dbi <= 8'h00;
		14'h3460:	ff_dbi <= 8'h00;
		14'h3461:	ff_dbi <= 8'h00;
		14'h3462:	ff_dbi <= 8'h00;
		14'h3463:	ff_dbi <= 8'h00;
		14'h3464:	ff_dbi <= 8'h00;
		14'h3465:	ff_dbi <= 8'h00;
		14'h3466:	ff_dbi <= 8'h00;
		14'h3467:	ff_dbi <= 8'h00;
		14'h3468:	ff_dbi <= 8'h00;
		14'h3469:	ff_dbi <= 8'h00;
		14'h346a:	ff_dbi <= 8'h00;
		14'h346b:	ff_dbi <= 8'h00;
		14'h346c:	ff_dbi <= 8'h00;
		14'h346d:	ff_dbi <= 8'h00;
		14'h346e:	ff_dbi <= 8'h00;
		14'h346f:	ff_dbi <= 8'h00;
		14'h3470:	ff_dbi <= 8'h00;
		14'h3471:	ff_dbi <= 8'h00;
		14'h3472:	ff_dbi <= 8'h00;
		14'h3473:	ff_dbi <= 8'h00;
		14'h3474:	ff_dbi <= 8'h00;
		14'h3475:	ff_dbi <= 8'h00;
		14'h3476:	ff_dbi <= 8'h00;
		14'h3477:	ff_dbi <= 8'h00;
		14'h3478:	ff_dbi <= 8'h00;
		14'h3479:	ff_dbi <= 8'h00;
		14'h347a:	ff_dbi <= 8'h00;
		14'h347b:	ff_dbi <= 8'h00;
		14'h347c:	ff_dbi <= 8'h00;
		14'h347d:	ff_dbi <= 8'h00;
		14'h347e:	ff_dbi <= 8'h00;
		14'h347f:	ff_dbi <= 8'h00;
		14'h3480:	ff_dbi <= 8'h00;
		14'h3481:	ff_dbi <= 8'h00;
		14'h3482:	ff_dbi <= 8'h00;
		14'h3483:	ff_dbi <= 8'h00;
		14'h3484:	ff_dbi <= 8'h00;
		14'h3485:	ff_dbi <= 8'h00;
		14'h3486:	ff_dbi <= 8'h00;
		14'h3487:	ff_dbi <= 8'h00;
		14'h3488:	ff_dbi <= 8'h00;
		14'h3489:	ff_dbi <= 8'h00;
		14'h348a:	ff_dbi <= 8'h00;
		14'h348b:	ff_dbi <= 8'h00;
		14'h348c:	ff_dbi <= 8'h00;
		14'h348d:	ff_dbi <= 8'h00;
		14'h348e:	ff_dbi <= 8'h00;
		14'h348f:	ff_dbi <= 8'h00;
		14'h3490:	ff_dbi <= 8'h00;
		14'h3491:	ff_dbi <= 8'h00;
		14'h3492:	ff_dbi <= 8'h00;
		14'h3493:	ff_dbi <= 8'h00;
		14'h3494:	ff_dbi <= 8'h00;
		14'h3495:	ff_dbi <= 8'h00;
		14'h3496:	ff_dbi <= 8'h00;
		14'h3497:	ff_dbi <= 8'h00;
		14'h3498:	ff_dbi <= 8'h00;
		14'h3499:	ff_dbi <= 8'h00;
		14'h349a:	ff_dbi <= 8'h00;
		14'h349b:	ff_dbi <= 8'h00;
		14'h349c:	ff_dbi <= 8'h00;
		14'h349d:	ff_dbi <= 8'h00;
		14'h349e:	ff_dbi <= 8'h00;
		14'h349f:	ff_dbi <= 8'h00;
		14'h34a0:	ff_dbi <= 8'h00;
		14'h34a1:	ff_dbi <= 8'h00;
		14'h34a2:	ff_dbi <= 8'h00;
		14'h34a3:	ff_dbi <= 8'h00;
		14'h34a4:	ff_dbi <= 8'h00;
		14'h34a5:	ff_dbi <= 8'h00;
		14'h34a6:	ff_dbi <= 8'h00;
		14'h34a7:	ff_dbi <= 8'h00;
		14'h34a8:	ff_dbi <= 8'h00;
		14'h34a9:	ff_dbi <= 8'h00;
		14'h34aa:	ff_dbi <= 8'h00;
		14'h34ab:	ff_dbi <= 8'h00;
		14'h34ac:	ff_dbi <= 8'h00;
		14'h34ad:	ff_dbi <= 8'h00;
		14'h34ae:	ff_dbi <= 8'h00;
		14'h34af:	ff_dbi <= 8'h00;
		14'h34b0:	ff_dbi <= 8'h00;
		14'h34b1:	ff_dbi <= 8'h00;
		14'h34b2:	ff_dbi <= 8'h00;
		14'h34b3:	ff_dbi <= 8'h00;
		14'h34b4:	ff_dbi <= 8'h00;
		14'h34b5:	ff_dbi <= 8'h00;
		14'h34b6:	ff_dbi <= 8'h00;
		14'h34b7:	ff_dbi <= 8'h00;
		14'h34b8:	ff_dbi <= 8'h00;
		14'h34b9:	ff_dbi <= 8'h00;
		14'h34ba:	ff_dbi <= 8'h00;
		14'h34bb:	ff_dbi <= 8'h00;
		14'h34bc:	ff_dbi <= 8'h00;
		14'h34bd:	ff_dbi <= 8'h00;
		14'h34be:	ff_dbi <= 8'h00;
		14'h34bf:	ff_dbi <= 8'h00;
		14'h34c0:	ff_dbi <= 8'h00;
		14'h34c1:	ff_dbi <= 8'h00;
		14'h34c2:	ff_dbi <= 8'h00;
		14'h34c3:	ff_dbi <= 8'h00;
		14'h34c4:	ff_dbi <= 8'h00;
		14'h34c5:	ff_dbi <= 8'h00;
		14'h34c6:	ff_dbi <= 8'h00;
		14'h34c7:	ff_dbi <= 8'h00;
		14'h34c8:	ff_dbi <= 8'h00;
		14'h34c9:	ff_dbi <= 8'h00;
		14'h34ca:	ff_dbi <= 8'h00;
		14'h34cb:	ff_dbi <= 8'h00;
		14'h34cc:	ff_dbi <= 8'h00;
		14'h34cd:	ff_dbi <= 8'h00;
		14'h34ce:	ff_dbi <= 8'h00;
		14'h34cf:	ff_dbi <= 8'h00;
		14'h34d0:	ff_dbi <= 8'h00;
		14'h34d1:	ff_dbi <= 8'h00;
		14'h34d2:	ff_dbi <= 8'h00;
		14'h34d3:	ff_dbi <= 8'h00;
		14'h34d4:	ff_dbi <= 8'h00;
		14'h34d5:	ff_dbi <= 8'h00;
		14'h34d6:	ff_dbi <= 8'h00;
		14'h34d7:	ff_dbi <= 8'h00;
		14'h34d8:	ff_dbi <= 8'h00;
		14'h34d9:	ff_dbi <= 8'h00;
		14'h34da:	ff_dbi <= 8'h00;
		14'h34db:	ff_dbi <= 8'h00;
		14'h34dc:	ff_dbi <= 8'h00;
		14'h34dd:	ff_dbi <= 8'h00;
		14'h34de:	ff_dbi <= 8'h00;
		14'h34df:	ff_dbi <= 8'h00;
		14'h34e0:	ff_dbi <= 8'h00;
		14'h34e1:	ff_dbi <= 8'h00;
		14'h34e2:	ff_dbi <= 8'h00;
		14'h34e3:	ff_dbi <= 8'h00;
		14'h34e4:	ff_dbi <= 8'h00;
		14'h34e5:	ff_dbi <= 8'h00;
		14'h34e6:	ff_dbi <= 8'h00;
		14'h34e7:	ff_dbi <= 8'h00;
		14'h34e8:	ff_dbi <= 8'h00;
		14'h34e9:	ff_dbi <= 8'h00;
		14'h34ea:	ff_dbi <= 8'h00;
		14'h34eb:	ff_dbi <= 8'h00;
		14'h34ec:	ff_dbi <= 8'h00;
		14'h34ed:	ff_dbi <= 8'h00;
		14'h34ee:	ff_dbi <= 8'h00;
		14'h34ef:	ff_dbi <= 8'h00;
		14'h34f0:	ff_dbi <= 8'h00;
		14'h34f1:	ff_dbi <= 8'h00;
		14'h34f2:	ff_dbi <= 8'h00;
		14'h34f3:	ff_dbi <= 8'h00;
		14'h34f4:	ff_dbi <= 8'h00;
		14'h34f5:	ff_dbi <= 8'h00;
		14'h34f6:	ff_dbi <= 8'h00;
		14'h34f7:	ff_dbi <= 8'h00;
		14'h34f8:	ff_dbi <= 8'h00;
		14'h34f9:	ff_dbi <= 8'h00;
		14'h34fa:	ff_dbi <= 8'h00;
		14'h34fb:	ff_dbi <= 8'h00;
		14'h34fc:	ff_dbi <= 8'h00;
		14'h34fd:	ff_dbi <= 8'h00;
		14'h34fe:	ff_dbi <= 8'h00;
		14'h34ff:	ff_dbi <= 8'h00;
		14'h3500:	ff_dbi <= 8'h00;
		14'h3501:	ff_dbi <= 8'h00;
		14'h3502:	ff_dbi <= 8'h00;
		14'h3503:	ff_dbi <= 8'h00;
		14'h3504:	ff_dbi <= 8'h00;
		14'h3505:	ff_dbi <= 8'h00;
		14'h3506:	ff_dbi <= 8'h00;
		14'h3507:	ff_dbi <= 8'h00;
		14'h3508:	ff_dbi <= 8'h00;
		14'h3509:	ff_dbi <= 8'h00;
		14'h350a:	ff_dbi <= 8'h00;
		14'h350b:	ff_dbi <= 8'h00;
		14'h350c:	ff_dbi <= 8'h00;
		14'h350d:	ff_dbi <= 8'h00;
		14'h350e:	ff_dbi <= 8'h00;
		14'h350f:	ff_dbi <= 8'h00;
		14'h3510:	ff_dbi <= 8'h00;
		14'h3511:	ff_dbi <= 8'h00;
		14'h3512:	ff_dbi <= 8'h00;
		14'h3513:	ff_dbi <= 8'h00;
		14'h3514:	ff_dbi <= 8'h00;
		14'h3515:	ff_dbi <= 8'h00;
		14'h3516:	ff_dbi <= 8'h00;
		14'h3517:	ff_dbi <= 8'h00;
		14'h3518:	ff_dbi <= 8'h00;
		14'h3519:	ff_dbi <= 8'h00;
		14'h351a:	ff_dbi <= 8'h00;
		14'h351b:	ff_dbi <= 8'h00;
		14'h351c:	ff_dbi <= 8'h00;
		14'h351d:	ff_dbi <= 8'h00;
		14'h351e:	ff_dbi <= 8'h00;
		14'h351f:	ff_dbi <= 8'h00;
		14'h3520:	ff_dbi <= 8'h00;
		14'h3521:	ff_dbi <= 8'h00;
		14'h3522:	ff_dbi <= 8'h00;
		14'h3523:	ff_dbi <= 8'h00;
		14'h3524:	ff_dbi <= 8'h00;
		14'h3525:	ff_dbi <= 8'h00;
		14'h3526:	ff_dbi <= 8'h00;
		14'h3527:	ff_dbi <= 8'h00;
		14'h3528:	ff_dbi <= 8'h00;
		14'h3529:	ff_dbi <= 8'h00;
		14'h352a:	ff_dbi <= 8'h00;
		14'h352b:	ff_dbi <= 8'h00;
		14'h352c:	ff_dbi <= 8'h00;
		14'h352d:	ff_dbi <= 8'h00;
		14'h352e:	ff_dbi <= 8'h00;
		14'h352f:	ff_dbi <= 8'h00;
		14'h3530:	ff_dbi <= 8'h00;
		14'h3531:	ff_dbi <= 8'h00;
		14'h3532:	ff_dbi <= 8'h00;
		14'h3533:	ff_dbi <= 8'h00;
		14'h3534:	ff_dbi <= 8'h00;
		14'h3535:	ff_dbi <= 8'h00;
		14'h3536:	ff_dbi <= 8'h00;
		14'h3537:	ff_dbi <= 8'h00;
		14'h3538:	ff_dbi <= 8'h00;
		14'h3539:	ff_dbi <= 8'h00;
		14'h353a:	ff_dbi <= 8'h00;
		14'h353b:	ff_dbi <= 8'h00;
		14'h353c:	ff_dbi <= 8'h00;
		14'h353d:	ff_dbi <= 8'h00;
		14'h353e:	ff_dbi <= 8'h00;
		14'h353f:	ff_dbi <= 8'h00;
		14'h3540:	ff_dbi <= 8'h00;
		14'h3541:	ff_dbi <= 8'h00;
		14'h3542:	ff_dbi <= 8'h00;
		14'h3543:	ff_dbi <= 8'h00;
		14'h3544:	ff_dbi <= 8'h00;
		14'h3545:	ff_dbi <= 8'h00;
		14'h3546:	ff_dbi <= 8'h00;
		14'h3547:	ff_dbi <= 8'h00;
		14'h3548:	ff_dbi <= 8'h00;
		14'h3549:	ff_dbi <= 8'h00;
		14'h354a:	ff_dbi <= 8'h00;
		14'h354b:	ff_dbi <= 8'h00;
		14'h354c:	ff_dbi <= 8'h00;
		14'h354d:	ff_dbi <= 8'h00;
		14'h354e:	ff_dbi <= 8'h00;
		14'h354f:	ff_dbi <= 8'h00;
		14'h3550:	ff_dbi <= 8'h00;
		14'h3551:	ff_dbi <= 8'h00;
		14'h3552:	ff_dbi <= 8'h00;
		14'h3553:	ff_dbi <= 8'h00;
		14'h3554:	ff_dbi <= 8'h00;
		14'h3555:	ff_dbi <= 8'h00;
		14'h3556:	ff_dbi <= 8'h00;
		14'h3557:	ff_dbi <= 8'h00;
		14'h3558:	ff_dbi <= 8'h00;
		14'h3559:	ff_dbi <= 8'h00;
		14'h355a:	ff_dbi <= 8'h00;
		14'h355b:	ff_dbi <= 8'h00;
		14'h355c:	ff_dbi <= 8'h00;
		14'h355d:	ff_dbi <= 8'h00;
		14'h355e:	ff_dbi <= 8'h00;
		14'h355f:	ff_dbi <= 8'h00;
		14'h3560:	ff_dbi <= 8'h00;
		14'h3561:	ff_dbi <= 8'h00;
		14'h3562:	ff_dbi <= 8'h00;
		14'h3563:	ff_dbi <= 8'h00;
		14'h3564:	ff_dbi <= 8'h00;
		14'h3565:	ff_dbi <= 8'h00;
		14'h3566:	ff_dbi <= 8'h00;
		14'h3567:	ff_dbi <= 8'h00;
		14'h3568:	ff_dbi <= 8'h00;
		14'h3569:	ff_dbi <= 8'h00;
		14'h356a:	ff_dbi <= 8'h00;
		14'h356b:	ff_dbi <= 8'h00;
		14'h356c:	ff_dbi <= 8'h00;
		14'h356d:	ff_dbi <= 8'h00;
		14'h356e:	ff_dbi <= 8'h00;
		14'h356f:	ff_dbi <= 8'h00;
		14'h3570:	ff_dbi <= 8'h00;
		14'h3571:	ff_dbi <= 8'h00;
		14'h3572:	ff_dbi <= 8'h00;
		14'h3573:	ff_dbi <= 8'h00;
		14'h3574:	ff_dbi <= 8'h00;
		14'h3575:	ff_dbi <= 8'h00;
		14'h3576:	ff_dbi <= 8'h00;
		14'h3577:	ff_dbi <= 8'h00;
		14'h3578:	ff_dbi <= 8'h00;
		14'h3579:	ff_dbi <= 8'h00;
		14'h357a:	ff_dbi <= 8'h00;
		14'h357b:	ff_dbi <= 8'h00;
		14'h357c:	ff_dbi <= 8'h00;
		14'h357d:	ff_dbi <= 8'h00;
		14'h357e:	ff_dbi <= 8'h00;
		14'h357f:	ff_dbi <= 8'h00;
		14'h3580:	ff_dbi <= 8'h00;
		14'h3581:	ff_dbi <= 8'h00;
		14'h3582:	ff_dbi <= 8'h00;
		14'h3583:	ff_dbi <= 8'h00;
		14'h3584:	ff_dbi <= 8'h00;
		14'h3585:	ff_dbi <= 8'h00;
		14'h3586:	ff_dbi <= 8'h00;
		14'h3587:	ff_dbi <= 8'h00;
		14'h3588:	ff_dbi <= 8'h00;
		14'h3589:	ff_dbi <= 8'h00;
		14'h358a:	ff_dbi <= 8'h00;
		14'h358b:	ff_dbi <= 8'h00;
		14'h358c:	ff_dbi <= 8'h00;
		14'h358d:	ff_dbi <= 8'h00;
		14'h358e:	ff_dbi <= 8'h00;
		14'h358f:	ff_dbi <= 8'h00;
		14'h3590:	ff_dbi <= 8'h00;
		14'h3591:	ff_dbi <= 8'h00;
		14'h3592:	ff_dbi <= 8'h00;
		14'h3593:	ff_dbi <= 8'h00;
		14'h3594:	ff_dbi <= 8'h00;
		14'h3595:	ff_dbi <= 8'h00;
		14'h3596:	ff_dbi <= 8'h00;
		14'h3597:	ff_dbi <= 8'h00;
		14'h3598:	ff_dbi <= 8'h00;
		14'h3599:	ff_dbi <= 8'h00;
		14'h359a:	ff_dbi <= 8'h00;
		14'h359b:	ff_dbi <= 8'h00;
		14'h359c:	ff_dbi <= 8'h00;
		14'h359d:	ff_dbi <= 8'h00;
		14'h359e:	ff_dbi <= 8'h00;
		14'h359f:	ff_dbi <= 8'h00;
		14'h35a0:	ff_dbi <= 8'h00;
		14'h35a1:	ff_dbi <= 8'h00;
		14'h35a2:	ff_dbi <= 8'h00;
		14'h35a3:	ff_dbi <= 8'h00;
		14'h35a4:	ff_dbi <= 8'h00;
		14'h35a5:	ff_dbi <= 8'h00;
		14'h35a6:	ff_dbi <= 8'h00;
		14'h35a7:	ff_dbi <= 8'h00;
		14'h35a8:	ff_dbi <= 8'h00;
		14'h35a9:	ff_dbi <= 8'h00;
		14'h35aa:	ff_dbi <= 8'h00;
		14'h35ab:	ff_dbi <= 8'h00;
		14'h35ac:	ff_dbi <= 8'h00;
		14'h35ad:	ff_dbi <= 8'h00;
		14'h35ae:	ff_dbi <= 8'h00;
		14'h35af:	ff_dbi <= 8'h00;
		14'h35b0:	ff_dbi <= 8'h00;
		14'h35b1:	ff_dbi <= 8'h00;
		14'h35b2:	ff_dbi <= 8'h00;
		14'h35b3:	ff_dbi <= 8'h00;
		14'h35b4:	ff_dbi <= 8'h00;
		14'h35b5:	ff_dbi <= 8'h00;
		14'h35b6:	ff_dbi <= 8'h00;
		14'h35b7:	ff_dbi <= 8'h00;
		14'h35b8:	ff_dbi <= 8'h00;
		14'h35b9:	ff_dbi <= 8'h00;
		14'h35ba:	ff_dbi <= 8'h00;
		14'h35bb:	ff_dbi <= 8'h00;
		14'h35bc:	ff_dbi <= 8'h00;
		14'h35bd:	ff_dbi <= 8'h00;
		14'h35be:	ff_dbi <= 8'h00;
		14'h35bf:	ff_dbi <= 8'h00;
		14'h35c0:	ff_dbi <= 8'h00;
		14'h35c1:	ff_dbi <= 8'h00;
		14'h35c2:	ff_dbi <= 8'h00;
		14'h35c3:	ff_dbi <= 8'h00;
		14'h35c4:	ff_dbi <= 8'h00;
		14'h35c5:	ff_dbi <= 8'h00;
		14'h35c6:	ff_dbi <= 8'h00;
		14'h35c7:	ff_dbi <= 8'h00;
		14'h35c8:	ff_dbi <= 8'h00;
		14'h35c9:	ff_dbi <= 8'h00;
		14'h35ca:	ff_dbi <= 8'h00;
		14'h35cb:	ff_dbi <= 8'h00;
		14'h35cc:	ff_dbi <= 8'h00;
		14'h35cd:	ff_dbi <= 8'h00;
		14'h35ce:	ff_dbi <= 8'h00;
		14'h35cf:	ff_dbi <= 8'h00;
		14'h35d0:	ff_dbi <= 8'h00;
		14'h35d1:	ff_dbi <= 8'h00;
		14'h35d2:	ff_dbi <= 8'h00;
		14'h35d3:	ff_dbi <= 8'h00;
		14'h35d4:	ff_dbi <= 8'h00;
		14'h35d5:	ff_dbi <= 8'h00;
		14'h35d6:	ff_dbi <= 8'h00;
		14'h35d7:	ff_dbi <= 8'h00;
		14'h35d8:	ff_dbi <= 8'h00;
		14'h35d9:	ff_dbi <= 8'h00;
		14'h35da:	ff_dbi <= 8'h00;
		14'h35db:	ff_dbi <= 8'h00;
		14'h35dc:	ff_dbi <= 8'h00;
		14'h35dd:	ff_dbi <= 8'h00;
		14'h35de:	ff_dbi <= 8'h00;
		14'h35df:	ff_dbi <= 8'h00;
		14'h35e0:	ff_dbi <= 8'h00;
		14'h35e1:	ff_dbi <= 8'h00;
		14'h35e2:	ff_dbi <= 8'h00;
		14'h35e3:	ff_dbi <= 8'h00;
		14'h35e4:	ff_dbi <= 8'h00;
		14'h35e5:	ff_dbi <= 8'h00;
		14'h35e6:	ff_dbi <= 8'h00;
		14'h35e7:	ff_dbi <= 8'h00;
		14'h35e8:	ff_dbi <= 8'h00;
		14'h35e9:	ff_dbi <= 8'h00;
		14'h35ea:	ff_dbi <= 8'h00;
		14'h35eb:	ff_dbi <= 8'h00;
		14'h35ec:	ff_dbi <= 8'h00;
		14'h35ed:	ff_dbi <= 8'h00;
		14'h35ee:	ff_dbi <= 8'h00;
		14'h35ef:	ff_dbi <= 8'h00;
		14'h35f0:	ff_dbi <= 8'h00;
		14'h35f1:	ff_dbi <= 8'h00;
		14'h35f2:	ff_dbi <= 8'h00;
		14'h35f3:	ff_dbi <= 8'h00;
		14'h35f4:	ff_dbi <= 8'h00;
		14'h35f5:	ff_dbi <= 8'h00;
		14'h35f6:	ff_dbi <= 8'h00;
		14'h35f7:	ff_dbi <= 8'h00;
		14'h35f8:	ff_dbi <= 8'h00;
		14'h35f9:	ff_dbi <= 8'h00;
		14'h35fa:	ff_dbi <= 8'h00;
		14'h35fb:	ff_dbi <= 8'h00;
		14'h35fc:	ff_dbi <= 8'h00;
		14'h35fd:	ff_dbi <= 8'h00;
		14'h35fe:	ff_dbi <= 8'h00;
		14'h35ff:	ff_dbi <= 8'h00;
		14'h3600:	ff_dbi <= 8'h00;
		14'h3601:	ff_dbi <= 8'h00;
		14'h3602:	ff_dbi <= 8'h00;
		14'h3603:	ff_dbi <= 8'h00;
		14'h3604:	ff_dbi <= 8'h00;
		14'h3605:	ff_dbi <= 8'h00;
		14'h3606:	ff_dbi <= 8'h00;
		14'h3607:	ff_dbi <= 8'h00;
		14'h3608:	ff_dbi <= 8'h00;
		14'h3609:	ff_dbi <= 8'h00;
		14'h360a:	ff_dbi <= 8'h00;
		14'h360b:	ff_dbi <= 8'h00;
		14'h360c:	ff_dbi <= 8'h00;
		14'h360d:	ff_dbi <= 8'h00;
		14'h360e:	ff_dbi <= 8'h00;
		14'h360f:	ff_dbi <= 8'h00;
		14'h3610:	ff_dbi <= 8'h00;
		14'h3611:	ff_dbi <= 8'h00;
		14'h3612:	ff_dbi <= 8'h00;
		14'h3613:	ff_dbi <= 8'h00;
		14'h3614:	ff_dbi <= 8'h00;
		14'h3615:	ff_dbi <= 8'h00;
		14'h3616:	ff_dbi <= 8'h00;
		14'h3617:	ff_dbi <= 8'h00;
		14'h3618:	ff_dbi <= 8'h00;
		14'h3619:	ff_dbi <= 8'h00;
		14'h361a:	ff_dbi <= 8'h00;
		14'h361b:	ff_dbi <= 8'h00;
		14'h361c:	ff_dbi <= 8'h00;
		14'h361d:	ff_dbi <= 8'h00;
		14'h361e:	ff_dbi <= 8'h00;
		14'h361f:	ff_dbi <= 8'h00;
		14'h3620:	ff_dbi <= 8'h00;
		14'h3621:	ff_dbi <= 8'h00;
		14'h3622:	ff_dbi <= 8'h00;
		14'h3623:	ff_dbi <= 8'h00;
		14'h3624:	ff_dbi <= 8'h00;
		14'h3625:	ff_dbi <= 8'h00;
		14'h3626:	ff_dbi <= 8'h00;
		14'h3627:	ff_dbi <= 8'h00;
		14'h3628:	ff_dbi <= 8'h00;
		14'h3629:	ff_dbi <= 8'h00;
		14'h362a:	ff_dbi <= 8'h00;
		14'h362b:	ff_dbi <= 8'h00;
		14'h362c:	ff_dbi <= 8'h00;
		14'h362d:	ff_dbi <= 8'h00;
		14'h362e:	ff_dbi <= 8'h00;
		14'h362f:	ff_dbi <= 8'h00;
		14'h3630:	ff_dbi <= 8'h00;
		14'h3631:	ff_dbi <= 8'h00;
		14'h3632:	ff_dbi <= 8'h00;
		14'h3633:	ff_dbi <= 8'h00;
		14'h3634:	ff_dbi <= 8'h00;
		14'h3635:	ff_dbi <= 8'h00;
		14'h3636:	ff_dbi <= 8'h00;
		14'h3637:	ff_dbi <= 8'h00;
		14'h3638:	ff_dbi <= 8'h00;
		14'h3639:	ff_dbi <= 8'h00;
		14'h363a:	ff_dbi <= 8'h00;
		14'h363b:	ff_dbi <= 8'h00;
		14'h363c:	ff_dbi <= 8'h00;
		14'h363d:	ff_dbi <= 8'h00;
		14'h363e:	ff_dbi <= 8'h00;
		14'h363f:	ff_dbi <= 8'h00;
		14'h3640:	ff_dbi <= 8'h00;
		14'h3641:	ff_dbi <= 8'h00;
		14'h3642:	ff_dbi <= 8'h00;
		14'h3643:	ff_dbi <= 8'h00;
		14'h3644:	ff_dbi <= 8'h00;
		14'h3645:	ff_dbi <= 8'h00;
		14'h3646:	ff_dbi <= 8'h00;
		14'h3647:	ff_dbi <= 8'h00;
		14'h3648:	ff_dbi <= 8'h00;
		14'h3649:	ff_dbi <= 8'h00;
		14'h364a:	ff_dbi <= 8'h00;
		14'h364b:	ff_dbi <= 8'h00;
		14'h364c:	ff_dbi <= 8'h00;
		14'h364d:	ff_dbi <= 8'h00;
		14'h364e:	ff_dbi <= 8'h00;
		14'h364f:	ff_dbi <= 8'h00;
		14'h3650:	ff_dbi <= 8'h00;
		14'h3651:	ff_dbi <= 8'h00;
		14'h3652:	ff_dbi <= 8'h00;
		14'h3653:	ff_dbi <= 8'h00;
		14'h3654:	ff_dbi <= 8'h00;
		14'h3655:	ff_dbi <= 8'h00;
		14'h3656:	ff_dbi <= 8'h00;
		14'h3657:	ff_dbi <= 8'h00;
		14'h3658:	ff_dbi <= 8'h00;
		14'h3659:	ff_dbi <= 8'h00;
		14'h365a:	ff_dbi <= 8'h00;
		14'h365b:	ff_dbi <= 8'h00;
		14'h365c:	ff_dbi <= 8'h00;
		14'h365d:	ff_dbi <= 8'h00;
		14'h365e:	ff_dbi <= 8'h00;
		14'h365f:	ff_dbi <= 8'h00;
		14'h3660:	ff_dbi <= 8'h00;
		14'h3661:	ff_dbi <= 8'h00;
		14'h3662:	ff_dbi <= 8'h00;
		14'h3663:	ff_dbi <= 8'h00;
		14'h3664:	ff_dbi <= 8'h00;
		14'h3665:	ff_dbi <= 8'h00;
		14'h3666:	ff_dbi <= 8'h00;
		14'h3667:	ff_dbi <= 8'h00;
		14'h3668:	ff_dbi <= 8'h00;
		14'h3669:	ff_dbi <= 8'h00;
		14'h366a:	ff_dbi <= 8'h00;
		14'h366b:	ff_dbi <= 8'h00;
		14'h366c:	ff_dbi <= 8'h00;
		14'h366d:	ff_dbi <= 8'h00;
		14'h366e:	ff_dbi <= 8'h00;
		14'h366f:	ff_dbi <= 8'h00;
		14'h3670:	ff_dbi <= 8'h00;
		14'h3671:	ff_dbi <= 8'h00;
		14'h3672:	ff_dbi <= 8'h00;
		14'h3673:	ff_dbi <= 8'h00;
		14'h3674:	ff_dbi <= 8'h00;
		14'h3675:	ff_dbi <= 8'h00;
		14'h3676:	ff_dbi <= 8'h00;
		14'h3677:	ff_dbi <= 8'h00;
		14'h3678:	ff_dbi <= 8'h00;
		14'h3679:	ff_dbi <= 8'h00;
		14'h367a:	ff_dbi <= 8'h00;
		14'h367b:	ff_dbi <= 8'h00;
		14'h367c:	ff_dbi <= 8'h00;
		14'h367d:	ff_dbi <= 8'h00;
		14'h367e:	ff_dbi <= 8'h00;
		14'h367f:	ff_dbi <= 8'h00;
		14'h3680:	ff_dbi <= 8'h00;
		14'h3681:	ff_dbi <= 8'h00;
		14'h3682:	ff_dbi <= 8'h00;
		14'h3683:	ff_dbi <= 8'h00;
		14'h3684:	ff_dbi <= 8'h00;
		14'h3685:	ff_dbi <= 8'h00;
		14'h3686:	ff_dbi <= 8'h00;
		14'h3687:	ff_dbi <= 8'h00;
		14'h3688:	ff_dbi <= 8'h00;
		14'h3689:	ff_dbi <= 8'h00;
		14'h368a:	ff_dbi <= 8'h00;
		14'h368b:	ff_dbi <= 8'h00;
		14'h368c:	ff_dbi <= 8'h00;
		14'h368d:	ff_dbi <= 8'h00;
		14'h368e:	ff_dbi <= 8'h00;
		14'h368f:	ff_dbi <= 8'h00;
		14'h3690:	ff_dbi <= 8'h00;
		14'h3691:	ff_dbi <= 8'h00;
		14'h3692:	ff_dbi <= 8'h00;
		14'h3693:	ff_dbi <= 8'h00;
		14'h3694:	ff_dbi <= 8'h00;
		14'h3695:	ff_dbi <= 8'h00;
		14'h3696:	ff_dbi <= 8'h00;
		14'h3697:	ff_dbi <= 8'h00;
		14'h3698:	ff_dbi <= 8'h00;
		14'h3699:	ff_dbi <= 8'h00;
		14'h369a:	ff_dbi <= 8'h00;
		14'h369b:	ff_dbi <= 8'h00;
		14'h369c:	ff_dbi <= 8'h00;
		14'h369d:	ff_dbi <= 8'h00;
		14'h369e:	ff_dbi <= 8'h00;
		14'h369f:	ff_dbi <= 8'h00;
		14'h36a0:	ff_dbi <= 8'h00;
		14'h36a1:	ff_dbi <= 8'h00;
		14'h36a2:	ff_dbi <= 8'h00;
		14'h36a3:	ff_dbi <= 8'h00;
		14'h36a4:	ff_dbi <= 8'h00;
		14'h36a5:	ff_dbi <= 8'h00;
		14'h36a6:	ff_dbi <= 8'h00;
		14'h36a7:	ff_dbi <= 8'h00;
		14'h36a8:	ff_dbi <= 8'h00;
		14'h36a9:	ff_dbi <= 8'h00;
		14'h36aa:	ff_dbi <= 8'h00;
		14'h36ab:	ff_dbi <= 8'h00;
		14'h36ac:	ff_dbi <= 8'h00;
		14'h36ad:	ff_dbi <= 8'h00;
		14'h36ae:	ff_dbi <= 8'h00;
		14'h36af:	ff_dbi <= 8'h00;
		14'h36b0:	ff_dbi <= 8'h00;
		14'h36b1:	ff_dbi <= 8'h00;
		14'h36b2:	ff_dbi <= 8'h00;
		14'h36b3:	ff_dbi <= 8'h00;
		14'h36b4:	ff_dbi <= 8'h00;
		14'h36b5:	ff_dbi <= 8'h00;
		14'h36b6:	ff_dbi <= 8'h00;
		14'h36b7:	ff_dbi <= 8'h00;
		14'h36b8:	ff_dbi <= 8'h00;
		14'h36b9:	ff_dbi <= 8'h00;
		14'h36ba:	ff_dbi <= 8'h00;
		14'h36bb:	ff_dbi <= 8'h00;
		14'h36bc:	ff_dbi <= 8'h00;
		14'h36bd:	ff_dbi <= 8'h00;
		14'h36be:	ff_dbi <= 8'h00;
		14'h36bf:	ff_dbi <= 8'h00;
		14'h36c0:	ff_dbi <= 8'h00;
		14'h36c1:	ff_dbi <= 8'h00;
		14'h36c2:	ff_dbi <= 8'h00;
		14'h36c3:	ff_dbi <= 8'h00;
		14'h36c4:	ff_dbi <= 8'h00;
		14'h36c5:	ff_dbi <= 8'h00;
		14'h36c6:	ff_dbi <= 8'h00;
		14'h36c7:	ff_dbi <= 8'h00;
		14'h36c8:	ff_dbi <= 8'h00;
		14'h36c9:	ff_dbi <= 8'h00;
		14'h36ca:	ff_dbi <= 8'h00;
		14'h36cb:	ff_dbi <= 8'h00;
		14'h36cc:	ff_dbi <= 8'h00;
		14'h36cd:	ff_dbi <= 8'h00;
		14'h36ce:	ff_dbi <= 8'h00;
		14'h36cf:	ff_dbi <= 8'h00;
		14'h36d0:	ff_dbi <= 8'h00;
		14'h36d1:	ff_dbi <= 8'h00;
		14'h36d2:	ff_dbi <= 8'h00;
		14'h36d3:	ff_dbi <= 8'h00;
		14'h36d4:	ff_dbi <= 8'h00;
		14'h36d5:	ff_dbi <= 8'h00;
		14'h36d6:	ff_dbi <= 8'h00;
		14'h36d7:	ff_dbi <= 8'h00;
		14'h36d8:	ff_dbi <= 8'h00;
		14'h36d9:	ff_dbi <= 8'h00;
		14'h36da:	ff_dbi <= 8'h00;
		14'h36db:	ff_dbi <= 8'h00;
		14'h36dc:	ff_dbi <= 8'h00;
		14'h36dd:	ff_dbi <= 8'h00;
		14'h36de:	ff_dbi <= 8'h00;
		14'h36df:	ff_dbi <= 8'h00;
		14'h36e0:	ff_dbi <= 8'h00;
		14'h36e1:	ff_dbi <= 8'h00;
		14'h36e2:	ff_dbi <= 8'h00;
		14'h36e3:	ff_dbi <= 8'h00;
		14'h36e4:	ff_dbi <= 8'h00;
		14'h36e5:	ff_dbi <= 8'h00;
		14'h36e6:	ff_dbi <= 8'h00;
		14'h36e7:	ff_dbi <= 8'h00;
		14'h36e8:	ff_dbi <= 8'h00;
		14'h36e9:	ff_dbi <= 8'h00;
		14'h36ea:	ff_dbi <= 8'h00;
		14'h36eb:	ff_dbi <= 8'h00;
		14'h36ec:	ff_dbi <= 8'h00;
		14'h36ed:	ff_dbi <= 8'h00;
		14'h36ee:	ff_dbi <= 8'h00;
		14'h36ef:	ff_dbi <= 8'h00;
		14'h36f0:	ff_dbi <= 8'h00;
		14'h36f1:	ff_dbi <= 8'h00;
		14'h36f2:	ff_dbi <= 8'h00;
		14'h36f3:	ff_dbi <= 8'h00;
		14'h36f4:	ff_dbi <= 8'h00;
		14'h36f5:	ff_dbi <= 8'h00;
		14'h36f6:	ff_dbi <= 8'h00;
		14'h36f7:	ff_dbi <= 8'h00;
		14'h36f8:	ff_dbi <= 8'h00;
		14'h36f9:	ff_dbi <= 8'h00;
		14'h36fa:	ff_dbi <= 8'h00;
		14'h36fb:	ff_dbi <= 8'h00;
		14'h36fc:	ff_dbi <= 8'h00;
		14'h36fd:	ff_dbi <= 8'h00;
		14'h36fe:	ff_dbi <= 8'h00;
		14'h36ff:	ff_dbi <= 8'h00;
		14'h3700:	ff_dbi <= 8'h00;
		14'h3701:	ff_dbi <= 8'h00;
		14'h3702:	ff_dbi <= 8'h00;
		14'h3703:	ff_dbi <= 8'h00;
		14'h3704:	ff_dbi <= 8'h00;
		14'h3705:	ff_dbi <= 8'h00;
		14'h3706:	ff_dbi <= 8'h00;
		14'h3707:	ff_dbi <= 8'h00;
		14'h3708:	ff_dbi <= 8'h00;
		14'h3709:	ff_dbi <= 8'h00;
		14'h370a:	ff_dbi <= 8'h00;
		14'h370b:	ff_dbi <= 8'h00;
		14'h370c:	ff_dbi <= 8'h00;
		14'h370d:	ff_dbi <= 8'h00;
		14'h370e:	ff_dbi <= 8'h00;
		14'h370f:	ff_dbi <= 8'h00;
		14'h3710:	ff_dbi <= 8'h00;
		14'h3711:	ff_dbi <= 8'h00;
		14'h3712:	ff_dbi <= 8'h00;
		14'h3713:	ff_dbi <= 8'h00;
		14'h3714:	ff_dbi <= 8'h00;
		14'h3715:	ff_dbi <= 8'h00;
		14'h3716:	ff_dbi <= 8'h00;
		14'h3717:	ff_dbi <= 8'h00;
		14'h3718:	ff_dbi <= 8'h00;
		14'h3719:	ff_dbi <= 8'h00;
		14'h371a:	ff_dbi <= 8'h00;
		14'h371b:	ff_dbi <= 8'h00;
		14'h371c:	ff_dbi <= 8'h00;
		14'h371d:	ff_dbi <= 8'h00;
		14'h371e:	ff_dbi <= 8'h00;
		14'h371f:	ff_dbi <= 8'h00;
		14'h3720:	ff_dbi <= 8'h00;
		14'h3721:	ff_dbi <= 8'h00;
		14'h3722:	ff_dbi <= 8'h00;
		14'h3723:	ff_dbi <= 8'h00;
		14'h3724:	ff_dbi <= 8'h00;
		14'h3725:	ff_dbi <= 8'h00;
		14'h3726:	ff_dbi <= 8'h00;
		14'h3727:	ff_dbi <= 8'h00;
		14'h3728:	ff_dbi <= 8'h00;
		14'h3729:	ff_dbi <= 8'h00;
		14'h372a:	ff_dbi <= 8'h00;
		14'h372b:	ff_dbi <= 8'h00;
		14'h372c:	ff_dbi <= 8'h00;
		14'h372d:	ff_dbi <= 8'h00;
		14'h372e:	ff_dbi <= 8'h00;
		14'h372f:	ff_dbi <= 8'h00;
		14'h3730:	ff_dbi <= 8'h00;
		14'h3731:	ff_dbi <= 8'h00;
		14'h3732:	ff_dbi <= 8'h00;
		14'h3733:	ff_dbi <= 8'h00;
		14'h3734:	ff_dbi <= 8'h00;
		14'h3735:	ff_dbi <= 8'h00;
		14'h3736:	ff_dbi <= 8'h00;
		14'h3737:	ff_dbi <= 8'h00;
		14'h3738:	ff_dbi <= 8'h00;
		14'h3739:	ff_dbi <= 8'h00;
		14'h373a:	ff_dbi <= 8'h00;
		14'h373b:	ff_dbi <= 8'h00;
		14'h373c:	ff_dbi <= 8'h00;
		14'h373d:	ff_dbi <= 8'h00;
		14'h373e:	ff_dbi <= 8'h00;
		14'h373f:	ff_dbi <= 8'h00;
		14'h3740:	ff_dbi <= 8'h00;
		14'h3741:	ff_dbi <= 8'h00;
		14'h3742:	ff_dbi <= 8'h00;
		14'h3743:	ff_dbi <= 8'h00;
		14'h3744:	ff_dbi <= 8'h00;
		14'h3745:	ff_dbi <= 8'h00;
		14'h3746:	ff_dbi <= 8'h00;
		14'h3747:	ff_dbi <= 8'h00;
		14'h3748:	ff_dbi <= 8'h00;
		14'h3749:	ff_dbi <= 8'h00;
		14'h374a:	ff_dbi <= 8'h00;
		14'h374b:	ff_dbi <= 8'h00;
		14'h374c:	ff_dbi <= 8'h00;
		14'h374d:	ff_dbi <= 8'h00;
		14'h374e:	ff_dbi <= 8'h00;
		14'h374f:	ff_dbi <= 8'h00;
		14'h3750:	ff_dbi <= 8'h00;
		14'h3751:	ff_dbi <= 8'h00;
		14'h3752:	ff_dbi <= 8'h00;
		14'h3753:	ff_dbi <= 8'h00;
		14'h3754:	ff_dbi <= 8'h00;
		14'h3755:	ff_dbi <= 8'h00;
		14'h3756:	ff_dbi <= 8'h00;
		14'h3757:	ff_dbi <= 8'h00;
		14'h3758:	ff_dbi <= 8'h00;
		14'h3759:	ff_dbi <= 8'h00;
		14'h375a:	ff_dbi <= 8'h00;
		14'h375b:	ff_dbi <= 8'h00;
		14'h375c:	ff_dbi <= 8'h00;
		14'h375d:	ff_dbi <= 8'h00;
		14'h375e:	ff_dbi <= 8'h00;
		14'h375f:	ff_dbi <= 8'h00;
		14'h3760:	ff_dbi <= 8'h00;
		14'h3761:	ff_dbi <= 8'h00;
		14'h3762:	ff_dbi <= 8'h00;
		14'h3763:	ff_dbi <= 8'h00;
		14'h3764:	ff_dbi <= 8'h00;
		14'h3765:	ff_dbi <= 8'h00;
		14'h3766:	ff_dbi <= 8'h00;
		14'h3767:	ff_dbi <= 8'h00;
		14'h3768:	ff_dbi <= 8'h00;
		14'h3769:	ff_dbi <= 8'h00;
		14'h376a:	ff_dbi <= 8'h00;
		14'h376b:	ff_dbi <= 8'h00;
		14'h376c:	ff_dbi <= 8'h00;
		14'h376d:	ff_dbi <= 8'h00;
		14'h376e:	ff_dbi <= 8'h00;
		14'h376f:	ff_dbi <= 8'h00;
		14'h3770:	ff_dbi <= 8'h00;
		14'h3771:	ff_dbi <= 8'h00;
		14'h3772:	ff_dbi <= 8'h00;
		14'h3773:	ff_dbi <= 8'h00;
		14'h3774:	ff_dbi <= 8'h00;
		14'h3775:	ff_dbi <= 8'h00;
		14'h3776:	ff_dbi <= 8'h00;
		14'h3777:	ff_dbi <= 8'h00;
		14'h3778:	ff_dbi <= 8'h00;
		14'h3779:	ff_dbi <= 8'h00;
		14'h377a:	ff_dbi <= 8'h00;
		14'h377b:	ff_dbi <= 8'h00;
		14'h377c:	ff_dbi <= 8'h00;
		14'h377d:	ff_dbi <= 8'h00;
		14'h377e:	ff_dbi <= 8'h00;
		14'h377f:	ff_dbi <= 8'h00;
		14'h3780:	ff_dbi <= 8'h00;
		14'h3781:	ff_dbi <= 8'h00;
		14'h3782:	ff_dbi <= 8'h00;
		14'h3783:	ff_dbi <= 8'h00;
		14'h3784:	ff_dbi <= 8'h00;
		14'h3785:	ff_dbi <= 8'h00;
		14'h3786:	ff_dbi <= 8'h00;
		14'h3787:	ff_dbi <= 8'h00;
		14'h3788:	ff_dbi <= 8'h00;
		14'h3789:	ff_dbi <= 8'h00;
		14'h378a:	ff_dbi <= 8'h00;
		14'h378b:	ff_dbi <= 8'h00;
		14'h378c:	ff_dbi <= 8'h00;
		14'h378d:	ff_dbi <= 8'h00;
		14'h378e:	ff_dbi <= 8'h00;
		14'h378f:	ff_dbi <= 8'h00;
		14'h3790:	ff_dbi <= 8'h00;
		14'h3791:	ff_dbi <= 8'h00;
		14'h3792:	ff_dbi <= 8'h00;
		14'h3793:	ff_dbi <= 8'h00;
		14'h3794:	ff_dbi <= 8'h00;
		14'h3795:	ff_dbi <= 8'h00;
		14'h3796:	ff_dbi <= 8'h00;
		14'h3797:	ff_dbi <= 8'h00;
		14'h3798:	ff_dbi <= 8'h00;
		14'h3799:	ff_dbi <= 8'h00;
		14'h379a:	ff_dbi <= 8'h00;
		14'h379b:	ff_dbi <= 8'h00;
		14'h379c:	ff_dbi <= 8'h00;
		14'h379d:	ff_dbi <= 8'h00;
		14'h379e:	ff_dbi <= 8'h00;
		14'h379f:	ff_dbi <= 8'h00;
		14'h37a0:	ff_dbi <= 8'h00;
		14'h37a1:	ff_dbi <= 8'h00;
		14'h37a2:	ff_dbi <= 8'h00;
		14'h37a3:	ff_dbi <= 8'h00;
		14'h37a4:	ff_dbi <= 8'h00;
		14'h37a5:	ff_dbi <= 8'h00;
		14'h37a6:	ff_dbi <= 8'h00;
		14'h37a7:	ff_dbi <= 8'h00;
		14'h37a8:	ff_dbi <= 8'h00;
		14'h37a9:	ff_dbi <= 8'h00;
		14'h37aa:	ff_dbi <= 8'h00;
		14'h37ab:	ff_dbi <= 8'h00;
		14'h37ac:	ff_dbi <= 8'h00;
		14'h37ad:	ff_dbi <= 8'h00;
		14'h37ae:	ff_dbi <= 8'h00;
		14'h37af:	ff_dbi <= 8'h00;
		14'h37b0:	ff_dbi <= 8'h00;
		14'h37b1:	ff_dbi <= 8'h00;
		14'h37b2:	ff_dbi <= 8'h00;
		14'h37b3:	ff_dbi <= 8'h00;
		14'h37b4:	ff_dbi <= 8'h00;
		14'h37b5:	ff_dbi <= 8'h00;
		14'h37b6:	ff_dbi <= 8'h00;
		14'h37b7:	ff_dbi <= 8'h00;
		14'h37b8:	ff_dbi <= 8'h00;
		14'h37b9:	ff_dbi <= 8'h00;
		14'h37ba:	ff_dbi <= 8'h00;
		14'h37bb:	ff_dbi <= 8'h00;
		14'h37bc:	ff_dbi <= 8'h00;
		14'h37bd:	ff_dbi <= 8'h00;
		14'h37be:	ff_dbi <= 8'h00;
		14'h37bf:	ff_dbi <= 8'h00;
		14'h37c0:	ff_dbi <= 8'h00;
		14'h37c1:	ff_dbi <= 8'h00;
		14'h37c2:	ff_dbi <= 8'h00;
		14'h37c3:	ff_dbi <= 8'h00;
		14'h37c4:	ff_dbi <= 8'h00;
		14'h37c5:	ff_dbi <= 8'h00;
		14'h37c6:	ff_dbi <= 8'h00;
		14'h37c7:	ff_dbi <= 8'h00;
		14'h37c8:	ff_dbi <= 8'h00;
		14'h37c9:	ff_dbi <= 8'h00;
		14'h37ca:	ff_dbi <= 8'h00;
		14'h37cb:	ff_dbi <= 8'h00;
		14'h37cc:	ff_dbi <= 8'h00;
		14'h37cd:	ff_dbi <= 8'h00;
		14'h37ce:	ff_dbi <= 8'h00;
		14'h37cf:	ff_dbi <= 8'h00;
		14'h37d0:	ff_dbi <= 8'h00;
		14'h37d1:	ff_dbi <= 8'h00;
		14'h37d2:	ff_dbi <= 8'h00;
		14'h37d3:	ff_dbi <= 8'h00;
		14'h37d4:	ff_dbi <= 8'h00;
		14'h37d5:	ff_dbi <= 8'h00;
		14'h37d6:	ff_dbi <= 8'h00;
		14'h37d7:	ff_dbi <= 8'h00;
		14'h37d8:	ff_dbi <= 8'h00;
		14'h37d9:	ff_dbi <= 8'h00;
		14'h37da:	ff_dbi <= 8'h00;
		14'h37db:	ff_dbi <= 8'h00;
		14'h37dc:	ff_dbi <= 8'h00;
		14'h37dd:	ff_dbi <= 8'h00;
		14'h37de:	ff_dbi <= 8'h00;
		14'h37df:	ff_dbi <= 8'h00;
		14'h37e0:	ff_dbi <= 8'h00;
		14'h37e1:	ff_dbi <= 8'h00;
		14'h37e2:	ff_dbi <= 8'h00;
		14'h37e3:	ff_dbi <= 8'h00;
		14'h37e4:	ff_dbi <= 8'h00;
		14'h37e5:	ff_dbi <= 8'h00;
		14'h37e6:	ff_dbi <= 8'h00;
		14'h37e7:	ff_dbi <= 8'h00;
		14'h37e8:	ff_dbi <= 8'h00;
		14'h37e9:	ff_dbi <= 8'h00;
		14'h37ea:	ff_dbi <= 8'h00;
		14'h37eb:	ff_dbi <= 8'h00;
		14'h37ec:	ff_dbi <= 8'h00;
		14'h37ed:	ff_dbi <= 8'h00;
		14'h37ee:	ff_dbi <= 8'h00;
		14'h37ef:	ff_dbi <= 8'h00;
		14'h37f0:	ff_dbi <= 8'h00;
		14'h37f1:	ff_dbi <= 8'h00;
		14'h37f2:	ff_dbi <= 8'h00;
		14'h37f3:	ff_dbi <= 8'h00;
		14'h37f4:	ff_dbi <= 8'h00;
		14'h37f5:	ff_dbi <= 8'h00;
		14'h37f6:	ff_dbi <= 8'h00;
		14'h37f7:	ff_dbi <= 8'h00;
		14'h37f8:	ff_dbi <= 8'h00;
		14'h37f9:	ff_dbi <= 8'h00;
		14'h37fa:	ff_dbi <= 8'h00;
		14'h37fb:	ff_dbi <= 8'h00;
		14'h37fc:	ff_dbi <= 8'h00;
		14'h37fd:	ff_dbi <= 8'h00;
		14'h37fe:	ff_dbi <= 8'h00;
		14'h37ff:	ff_dbi <= 8'h00;
		14'h3800:	ff_dbi <= 8'h00;
		14'h3801:	ff_dbi <= 8'h00;
		14'h3802:	ff_dbi <= 8'h00;
		14'h3803:	ff_dbi <= 8'h00;
		14'h3804:	ff_dbi <= 8'h00;
		14'h3805:	ff_dbi <= 8'h00;
		14'h3806:	ff_dbi <= 8'h00;
		14'h3807:	ff_dbi <= 8'h00;
		14'h3808:	ff_dbi <= 8'h00;
		14'h3809:	ff_dbi <= 8'h00;
		14'h380a:	ff_dbi <= 8'h00;
		14'h380b:	ff_dbi <= 8'h00;
		14'h380c:	ff_dbi <= 8'h00;
		14'h380d:	ff_dbi <= 8'h00;
		14'h380e:	ff_dbi <= 8'h00;
		14'h380f:	ff_dbi <= 8'h00;
		14'h3810:	ff_dbi <= 8'h00;
		14'h3811:	ff_dbi <= 8'h00;
		14'h3812:	ff_dbi <= 8'h00;
		14'h3813:	ff_dbi <= 8'h00;
		14'h3814:	ff_dbi <= 8'h00;
		14'h3815:	ff_dbi <= 8'h00;
		14'h3816:	ff_dbi <= 8'h00;
		14'h3817:	ff_dbi <= 8'h00;
		14'h3818:	ff_dbi <= 8'h00;
		14'h3819:	ff_dbi <= 8'h00;
		14'h381a:	ff_dbi <= 8'h00;
		14'h381b:	ff_dbi <= 8'h00;
		14'h381c:	ff_dbi <= 8'h00;
		14'h381d:	ff_dbi <= 8'h00;
		14'h381e:	ff_dbi <= 8'h00;
		14'h381f:	ff_dbi <= 8'h00;
		14'h3820:	ff_dbi <= 8'h00;
		14'h3821:	ff_dbi <= 8'h00;
		14'h3822:	ff_dbi <= 8'h00;
		14'h3823:	ff_dbi <= 8'h00;
		14'h3824:	ff_dbi <= 8'h00;
		14'h3825:	ff_dbi <= 8'h00;
		14'h3826:	ff_dbi <= 8'h00;
		14'h3827:	ff_dbi <= 8'h00;
		14'h3828:	ff_dbi <= 8'h00;
		14'h3829:	ff_dbi <= 8'h00;
		14'h382a:	ff_dbi <= 8'h00;
		14'h382b:	ff_dbi <= 8'h00;
		14'h382c:	ff_dbi <= 8'h00;
		14'h382d:	ff_dbi <= 8'h00;
		14'h382e:	ff_dbi <= 8'h00;
		14'h382f:	ff_dbi <= 8'h00;
		14'h3830:	ff_dbi <= 8'h00;
		14'h3831:	ff_dbi <= 8'h00;
		14'h3832:	ff_dbi <= 8'h00;
		14'h3833:	ff_dbi <= 8'h00;
		14'h3834:	ff_dbi <= 8'h00;
		14'h3835:	ff_dbi <= 8'h00;
		14'h3836:	ff_dbi <= 8'h00;
		14'h3837:	ff_dbi <= 8'h00;
		14'h3838:	ff_dbi <= 8'h00;
		14'h3839:	ff_dbi <= 8'h00;
		14'h383a:	ff_dbi <= 8'h00;
		14'h383b:	ff_dbi <= 8'h00;
		14'h383c:	ff_dbi <= 8'h00;
		14'h383d:	ff_dbi <= 8'h00;
		14'h383e:	ff_dbi <= 8'h00;
		14'h383f:	ff_dbi <= 8'h00;
		14'h3840:	ff_dbi <= 8'h00;
		14'h3841:	ff_dbi <= 8'h00;
		14'h3842:	ff_dbi <= 8'h00;
		14'h3843:	ff_dbi <= 8'h00;
		14'h3844:	ff_dbi <= 8'h00;
		14'h3845:	ff_dbi <= 8'h00;
		14'h3846:	ff_dbi <= 8'h00;
		14'h3847:	ff_dbi <= 8'h00;
		14'h3848:	ff_dbi <= 8'h00;
		14'h3849:	ff_dbi <= 8'h00;
		14'h384a:	ff_dbi <= 8'h00;
		14'h384b:	ff_dbi <= 8'h00;
		14'h384c:	ff_dbi <= 8'h00;
		14'h384d:	ff_dbi <= 8'h00;
		14'h384e:	ff_dbi <= 8'h00;
		14'h384f:	ff_dbi <= 8'h00;
		14'h3850:	ff_dbi <= 8'h00;
		14'h3851:	ff_dbi <= 8'h00;
		14'h3852:	ff_dbi <= 8'h00;
		14'h3853:	ff_dbi <= 8'h00;
		14'h3854:	ff_dbi <= 8'h00;
		14'h3855:	ff_dbi <= 8'h00;
		14'h3856:	ff_dbi <= 8'h00;
		14'h3857:	ff_dbi <= 8'h00;
		14'h3858:	ff_dbi <= 8'h00;
		14'h3859:	ff_dbi <= 8'h00;
		14'h385a:	ff_dbi <= 8'h00;
		14'h385b:	ff_dbi <= 8'h00;
		14'h385c:	ff_dbi <= 8'h00;
		14'h385d:	ff_dbi <= 8'h00;
		14'h385e:	ff_dbi <= 8'h00;
		14'h385f:	ff_dbi <= 8'h00;
		14'h3860:	ff_dbi <= 8'h00;
		14'h3861:	ff_dbi <= 8'h00;
		14'h3862:	ff_dbi <= 8'h00;
		14'h3863:	ff_dbi <= 8'h00;
		14'h3864:	ff_dbi <= 8'h00;
		14'h3865:	ff_dbi <= 8'h00;
		14'h3866:	ff_dbi <= 8'h00;
		14'h3867:	ff_dbi <= 8'h00;
		14'h3868:	ff_dbi <= 8'h00;
		14'h3869:	ff_dbi <= 8'h00;
		14'h386a:	ff_dbi <= 8'h00;
		14'h386b:	ff_dbi <= 8'h00;
		14'h386c:	ff_dbi <= 8'h00;
		14'h386d:	ff_dbi <= 8'h00;
		14'h386e:	ff_dbi <= 8'h00;
		14'h386f:	ff_dbi <= 8'h00;
		14'h3870:	ff_dbi <= 8'h00;
		14'h3871:	ff_dbi <= 8'h00;
		14'h3872:	ff_dbi <= 8'h00;
		14'h3873:	ff_dbi <= 8'h00;
		14'h3874:	ff_dbi <= 8'h00;
		14'h3875:	ff_dbi <= 8'h00;
		14'h3876:	ff_dbi <= 8'h00;
		14'h3877:	ff_dbi <= 8'h00;
		14'h3878:	ff_dbi <= 8'h00;
		14'h3879:	ff_dbi <= 8'h00;
		14'h387a:	ff_dbi <= 8'h00;
		14'h387b:	ff_dbi <= 8'h00;
		14'h387c:	ff_dbi <= 8'h00;
		14'h387d:	ff_dbi <= 8'h00;
		14'h387e:	ff_dbi <= 8'h00;
		14'h387f:	ff_dbi <= 8'h00;
		14'h3880:	ff_dbi <= 8'h00;
		14'h3881:	ff_dbi <= 8'h00;
		14'h3882:	ff_dbi <= 8'h00;
		14'h3883:	ff_dbi <= 8'h00;
		14'h3884:	ff_dbi <= 8'h00;
		14'h3885:	ff_dbi <= 8'h00;
		14'h3886:	ff_dbi <= 8'h00;
		14'h3887:	ff_dbi <= 8'h00;
		14'h3888:	ff_dbi <= 8'h00;
		14'h3889:	ff_dbi <= 8'h00;
		14'h388a:	ff_dbi <= 8'h00;
		14'h388b:	ff_dbi <= 8'h00;
		14'h388c:	ff_dbi <= 8'h00;
		14'h388d:	ff_dbi <= 8'h00;
		14'h388e:	ff_dbi <= 8'h00;
		14'h388f:	ff_dbi <= 8'h00;
		14'h3890:	ff_dbi <= 8'h00;
		14'h3891:	ff_dbi <= 8'h00;
		14'h3892:	ff_dbi <= 8'h00;
		14'h3893:	ff_dbi <= 8'h00;
		14'h3894:	ff_dbi <= 8'h00;
		14'h3895:	ff_dbi <= 8'h00;
		14'h3896:	ff_dbi <= 8'h00;
		14'h3897:	ff_dbi <= 8'h00;
		14'h3898:	ff_dbi <= 8'h00;
		14'h3899:	ff_dbi <= 8'h00;
		14'h389a:	ff_dbi <= 8'h00;
		14'h389b:	ff_dbi <= 8'h00;
		14'h389c:	ff_dbi <= 8'h00;
		14'h389d:	ff_dbi <= 8'h00;
		14'h389e:	ff_dbi <= 8'h00;
		14'h389f:	ff_dbi <= 8'h00;
		14'h38a0:	ff_dbi <= 8'h00;
		14'h38a1:	ff_dbi <= 8'h00;
		14'h38a2:	ff_dbi <= 8'h00;
		14'h38a3:	ff_dbi <= 8'h00;
		14'h38a4:	ff_dbi <= 8'h00;
		14'h38a5:	ff_dbi <= 8'h00;
		14'h38a6:	ff_dbi <= 8'h00;
		14'h38a7:	ff_dbi <= 8'h00;
		14'h38a8:	ff_dbi <= 8'h00;
		14'h38a9:	ff_dbi <= 8'h00;
		14'h38aa:	ff_dbi <= 8'h00;
		14'h38ab:	ff_dbi <= 8'h00;
		14'h38ac:	ff_dbi <= 8'h00;
		14'h38ad:	ff_dbi <= 8'h00;
		14'h38ae:	ff_dbi <= 8'h00;
		14'h38af:	ff_dbi <= 8'h00;
		14'h38b0:	ff_dbi <= 8'h00;
		14'h38b1:	ff_dbi <= 8'h00;
		14'h38b2:	ff_dbi <= 8'h00;
		14'h38b3:	ff_dbi <= 8'h00;
		14'h38b4:	ff_dbi <= 8'h00;
		14'h38b5:	ff_dbi <= 8'h00;
		14'h38b6:	ff_dbi <= 8'h00;
		14'h38b7:	ff_dbi <= 8'h00;
		14'h38b8:	ff_dbi <= 8'h00;
		14'h38b9:	ff_dbi <= 8'h00;
		14'h38ba:	ff_dbi <= 8'h00;
		14'h38bb:	ff_dbi <= 8'h00;
		14'h38bc:	ff_dbi <= 8'h00;
		14'h38bd:	ff_dbi <= 8'h00;
		14'h38be:	ff_dbi <= 8'h00;
		14'h38bf:	ff_dbi <= 8'h00;
		14'h38c0:	ff_dbi <= 8'h00;
		14'h38c1:	ff_dbi <= 8'h00;
		14'h38c2:	ff_dbi <= 8'h00;
		14'h38c3:	ff_dbi <= 8'h00;
		14'h38c4:	ff_dbi <= 8'h00;
		14'h38c5:	ff_dbi <= 8'h00;
		14'h38c6:	ff_dbi <= 8'h00;
		14'h38c7:	ff_dbi <= 8'h00;
		14'h38c8:	ff_dbi <= 8'h00;
		14'h38c9:	ff_dbi <= 8'h00;
		14'h38ca:	ff_dbi <= 8'h00;
		14'h38cb:	ff_dbi <= 8'h00;
		14'h38cc:	ff_dbi <= 8'h00;
		14'h38cd:	ff_dbi <= 8'h00;
		14'h38ce:	ff_dbi <= 8'h00;
		14'h38cf:	ff_dbi <= 8'h00;
		14'h38d0:	ff_dbi <= 8'h00;
		14'h38d1:	ff_dbi <= 8'h00;
		14'h38d2:	ff_dbi <= 8'h00;
		14'h38d3:	ff_dbi <= 8'h00;
		14'h38d4:	ff_dbi <= 8'h00;
		14'h38d5:	ff_dbi <= 8'h00;
		14'h38d6:	ff_dbi <= 8'h00;
		14'h38d7:	ff_dbi <= 8'h00;
		14'h38d8:	ff_dbi <= 8'h00;
		14'h38d9:	ff_dbi <= 8'h00;
		14'h38da:	ff_dbi <= 8'h00;
		14'h38db:	ff_dbi <= 8'h00;
		14'h38dc:	ff_dbi <= 8'h00;
		14'h38dd:	ff_dbi <= 8'h00;
		14'h38de:	ff_dbi <= 8'h00;
		14'h38df:	ff_dbi <= 8'h00;
		14'h38e0:	ff_dbi <= 8'h00;
		14'h38e1:	ff_dbi <= 8'h00;
		14'h38e2:	ff_dbi <= 8'h00;
		14'h38e3:	ff_dbi <= 8'h00;
		14'h38e4:	ff_dbi <= 8'h00;
		14'h38e5:	ff_dbi <= 8'h00;
		14'h38e6:	ff_dbi <= 8'h00;
		14'h38e7:	ff_dbi <= 8'h00;
		14'h38e8:	ff_dbi <= 8'h00;
		14'h38e9:	ff_dbi <= 8'h00;
		14'h38ea:	ff_dbi <= 8'h00;
		14'h38eb:	ff_dbi <= 8'h00;
		14'h38ec:	ff_dbi <= 8'h00;
		14'h38ed:	ff_dbi <= 8'h00;
		14'h38ee:	ff_dbi <= 8'h00;
		14'h38ef:	ff_dbi <= 8'h00;
		14'h38f0:	ff_dbi <= 8'h00;
		14'h38f1:	ff_dbi <= 8'h00;
		14'h38f2:	ff_dbi <= 8'h00;
		14'h38f3:	ff_dbi <= 8'h00;
		14'h38f4:	ff_dbi <= 8'h00;
		14'h38f5:	ff_dbi <= 8'h00;
		14'h38f6:	ff_dbi <= 8'h00;
		14'h38f7:	ff_dbi <= 8'h00;
		14'h38f8:	ff_dbi <= 8'h00;
		14'h38f9:	ff_dbi <= 8'h00;
		14'h38fa:	ff_dbi <= 8'h00;
		14'h38fb:	ff_dbi <= 8'h00;
		14'h38fc:	ff_dbi <= 8'h00;
		14'h38fd:	ff_dbi <= 8'h00;
		14'h38fe:	ff_dbi <= 8'h00;
		14'h38ff:	ff_dbi <= 8'h00;
		14'h3900:	ff_dbi <= 8'h00;
		14'h3901:	ff_dbi <= 8'h00;
		14'h3902:	ff_dbi <= 8'h00;
		14'h3903:	ff_dbi <= 8'h00;
		14'h3904:	ff_dbi <= 8'h00;
		14'h3905:	ff_dbi <= 8'h00;
		14'h3906:	ff_dbi <= 8'h00;
		14'h3907:	ff_dbi <= 8'h00;
		14'h3908:	ff_dbi <= 8'h00;
		14'h3909:	ff_dbi <= 8'h00;
		14'h390a:	ff_dbi <= 8'h00;
		14'h390b:	ff_dbi <= 8'h00;
		14'h390c:	ff_dbi <= 8'h00;
		14'h390d:	ff_dbi <= 8'h00;
		14'h390e:	ff_dbi <= 8'h00;
		14'h390f:	ff_dbi <= 8'h00;
		14'h3910:	ff_dbi <= 8'h00;
		14'h3911:	ff_dbi <= 8'h00;
		14'h3912:	ff_dbi <= 8'h00;
		14'h3913:	ff_dbi <= 8'h00;
		14'h3914:	ff_dbi <= 8'h00;
		14'h3915:	ff_dbi <= 8'h00;
		14'h3916:	ff_dbi <= 8'h00;
		14'h3917:	ff_dbi <= 8'h00;
		14'h3918:	ff_dbi <= 8'h00;
		14'h3919:	ff_dbi <= 8'h00;
		14'h391a:	ff_dbi <= 8'h00;
		14'h391b:	ff_dbi <= 8'h00;
		14'h391c:	ff_dbi <= 8'h00;
		14'h391d:	ff_dbi <= 8'h00;
		14'h391e:	ff_dbi <= 8'h00;
		14'h391f:	ff_dbi <= 8'h00;
		14'h3920:	ff_dbi <= 8'h00;
		14'h3921:	ff_dbi <= 8'h00;
		14'h3922:	ff_dbi <= 8'h00;
		14'h3923:	ff_dbi <= 8'h00;
		14'h3924:	ff_dbi <= 8'h00;
		14'h3925:	ff_dbi <= 8'h00;
		14'h3926:	ff_dbi <= 8'h00;
		14'h3927:	ff_dbi <= 8'h00;
		14'h3928:	ff_dbi <= 8'h00;
		14'h3929:	ff_dbi <= 8'h00;
		14'h392a:	ff_dbi <= 8'h00;
		14'h392b:	ff_dbi <= 8'h00;
		14'h392c:	ff_dbi <= 8'h00;
		14'h392d:	ff_dbi <= 8'h00;
		14'h392e:	ff_dbi <= 8'h00;
		14'h392f:	ff_dbi <= 8'h00;
		14'h3930:	ff_dbi <= 8'h00;
		14'h3931:	ff_dbi <= 8'h00;
		14'h3932:	ff_dbi <= 8'h00;
		14'h3933:	ff_dbi <= 8'h00;
		14'h3934:	ff_dbi <= 8'h00;
		14'h3935:	ff_dbi <= 8'h00;
		14'h3936:	ff_dbi <= 8'h00;
		14'h3937:	ff_dbi <= 8'h00;
		14'h3938:	ff_dbi <= 8'h00;
		14'h3939:	ff_dbi <= 8'h00;
		14'h393a:	ff_dbi <= 8'h00;
		14'h393b:	ff_dbi <= 8'h00;
		14'h393c:	ff_dbi <= 8'h00;
		14'h393d:	ff_dbi <= 8'h00;
		14'h393e:	ff_dbi <= 8'h00;
		14'h393f:	ff_dbi <= 8'h00;
		14'h3940:	ff_dbi <= 8'h00;
		14'h3941:	ff_dbi <= 8'h00;
		14'h3942:	ff_dbi <= 8'h00;
		14'h3943:	ff_dbi <= 8'h00;
		14'h3944:	ff_dbi <= 8'h00;
		14'h3945:	ff_dbi <= 8'h00;
		14'h3946:	ff_dbi <= 8'h00;
		14'h3947:	ff_dbi <= 8'h00;
		14'h3948:	ff_dbi <= 8'h00;
		14'h3949:	ff_dbi <= 8'h00;
		14'h394a:	ff_dbi <= 8'h00;
		14'h394b:	ff_dbi <= 8'h00;
		14'h394c:	ff_dbi <= 8'h00;
		14'h394d:	ff_dbi <= 8'h00;
		14'h394e:	ff_dbi <= 8'h00;
		14'h394f:	ff_dbi <= 8'h00;
		14'h3950:	ff_dbi <= 8'h00;
		14'h3951:	ff_dbi <= 8'h00;
		14'h3952:	ff_dbi <= 8'h00;
		14'h3953:	ff_dbi <= 8'h00;
		14'h3954:	ff_dbi <= 8'h00;
		14'h3955:	ff_dbi <= 8'h00;
		14'h3956:	ff_dbi <= 8'h00;
		14'h3957:	ff_dbi <= 8'h00;
		14'h3958:	ff_dbi <= 8'h00;
		14'h3959:	ff_dbi <= 8'h00;
		14'h395a:	ff_dbi <= 8'h00;
		14'h395b:	ff_dbi <= 8'h00;
		14'h395c:	ff_dbi <= 8'h00;
		14'h395d:	ff_dbi <= 8'h00;
		14'h395e:	ff_dbi <= 8'h00;
		14'h395f:	ff_dbi <= 8'h00;
		14'h3960:	ff_dbi <= 8'h00;
		14'h3961:	ff_dbi <= 8'h00;
		14'h3962:	ff_dbi <= 8'h00;
		14'h3963:	ff_dbi <= 8'h00;
		14'h3964:	ff_dbi <= 8'h00;
		14'h3965:	ff_dbi <= 8'h00;
		14'h3966:	ff_dbi <= 8'h00;
		14'h3967:	ff_dbi <= 8'h00;
		14'h3968:	ff_dbi <= 8'h00;
		14'h3969:	ff_dbi <= 8'h00;
		14'h396a:	ff_dbi <= 8'h00;
		14'h396b:	ff_dbi <= 8'h00;
		14'h396c:	ff_dbi <= 8'h00;
		14'h396d:	ff_dbi <= 8'h00;
		14'h396e:	ff_dbi <= 8'h00;
		14'h396f:	ff_dbi <= 8'h00;
		14'h3970:	ff_dbi <= 8'h00;
		14'h3971:	ff_dbi <= 8'h00;
		14'h3972:	ff_dbi <= 8'h00;
		14'h3973:	ff_dbi <= 8'h00;
		14'h3974:	ff_dbi <= 8'h00;
		14'h3975:	ff_dbi <= 8'h00;
		14'h3976:	ff_dbi <= 8'h00;
		14'h3977:	ff_dbi <= 8'h00;
		14'h3978:	ff_dbi <= 8'h00;
		14'h3979:	ff_dbi <= 8'h00;
		14'h397a:	ff_dbi <= 8'h00;
		14'h397b:	ff_dbi <= 8'h00;
		14'h397c:	ff_dbi <= 8'h00;
		14'h397d:	ff_dbi <= 8'h00;
		14'h397e:	ff_dbi <= 8'h00;
		14'h397f:	ff_dbi <= 8'h00;
		14'h3980:	ff_dbi <= 8'h00;
		14'h3981:	ff_dbi <= 8'h00;
		14'h3982:	ff_dbi <= 8'h00;
		14'h3983:	ff_dbi <= 8'h00;
		14'h3984:	ff_dbi <= 8'h00;
		14'h3985:	ff_dbi <= 8'h00;
		14'h3986:	ff_dbi <= 8'h00;
		14'h3987:	ff_dbi <= 8'h00;
		14'h3988:	ff_dbi <= 8'h00;
		14'h3989:	ff_dbi <= 8'h00;
		14'h398a:	ff_dbi <= 8'h00;
		14'h398b:	ff_dbi <= 8'h00;
		14'h398c:	ff_dbi <= 8'h00;
		14'h398d:	ff_dbi <= 8'h00;
		14'h398e:	ff_dbi <= 8'h00;
		14'h398f:	ff_dbi <= 8'h00;
		14'h3990:	ff_dbi <= 8'h00;
		14'h3991:	ff_dbi <= 8'h00;
		14'h3992:	ff_dbi <= 8'h00;
		14'h3993:	ff_dbi <= 8'h00;
		14'h3994:	ff_dbi <= 8'h00;
		14'h3995:	ff_dbi <= 8'h00;
		14'h3996:	ff_dbi <= 8'h00;
		14'h3997:	ff_dbi <= 8'h00;
		14'h3998:	ff_dbi <= 8'h00;
		14'h3999:	ff_dbi <= 8'h00;
		14'h399a:	ff_dbi <= 8'h00;
		14'h399b:	ff_dbi <= 8'h00;
		14'h399c:	ff_dbi <= 8'h00;
		14'h399d:	ff_dbi <= 8'h00;
		14'h399e:	ff_dbi <= 8'h00;
		14'h399f:	ff_dbi <= 8'h00;
		14'h39a0:	ff_dbi <= 8'h00;
		14'h39a1:	ff_dbi <= 8'h00;
		14'h39a2:	ff_dbi <= 8'h00;
		14'h39a3:	ff_dbi <= 8'h00;
		14'h39a4:	ff_dbi <= 8'h00;
		14'h39a5:	ff_dbi <= 8'h00;
		14'h39a6:	ff_dbi <= 8'h00;
		14'h39a7:	ff_dbi <= 8'h00;
		14'h39a8:	ff_dbi <= 8'h00;
		14'h39a9:	ff_dbi <= 8'h00;
		14'h39aa:	ff_dbi <= 8'h00;
		14'h39ab:	ff_dbi <= 8'h00;
		14'h39ac:	ff_dbi <= 8'h00;
		14'h39ad:	ff_dbi <= 8'h00;
		14'h39ae:	ff_dbi <= 8'h00;
		14'h39af:	ff_dbi <= 8'h00;
		14'h39b0:	ff_dbi <= 8'h00;
		14'h39b1:	ff_dbi <= 8'h00;
		14'h39b2:	ff_dbi <= 8'h00;
		14'h39b3:	ff_dbi <= 8'h00;
		14'h39b4:	ff_dbi <= 8'h00;
		14'h39b5:	ff_dbi <= 8'h00;
		14'h39b6:	ff_dbi <= 8'h00;
		14'h39b7:	ff_dbi <= 8'h00;
		14'h39b8:	ff_dbi <= 8'h00;
		14'h39b9:	ff_dbi <= 8'h00;
		14'h39ba:	ff_dbi <= 8'h00;
		14'h39bb:	ff_dbi <= 8'h00;
		14'h39bc:	ff_dbi <= 8'h00;
		14'h39bd:	ff_dbi <= 8'h00;
		14'h39be:	ff_dbi <= 8'h00;
		14'h39bf:	ff_dbi <= 8'h00;
		14'h39c0:	ff_dbi <= 8'h00;
		14'h39c1:	ff_dbi <= 8'h00;
		14'h39c2:	ff_dbi <= 8'h00;
		14'h39c3:	ff_dbi <= 8'h00;
		14'h39c4:	ff_dbi <= 8'h00;
		14'h39c5:	ff_dbi <= 8'h00;
		14'h39c6:	ff_dbi <= 8'h00;
		14'h39c7:	ff_dbi <= 8'h00;
		14'h39c8:	ff_dbi <= 8'h00;
		14'h39c9:	ff_dbi <= 8'h00;
		14'h39ca:	ff_dbi <= 8'h00;
		14'h39cb:	ff_dbi <= 8'h00;
		14'h39cc:	ff_dbi <= 8'h00;
		14'h39cd:	ff_dbi <= 8'h00;
		14'h39ce:	ff_dbi <= 8'h00;
		14'h39cf:	ff_dbi <= 8'h00;
		14'h39d0:	ff_dbi <= 8'h00;
		14'h39d1:	ff_dbi <= 8'h00;
		14'h39d2:	ff_dbi <= 8'h00;
		14'h39d3:	ff_dbi <= 8'h00;
		14'h39d4:	ff_dbi <= 8'h00;
		14'h39d5:	ff_dbi <= 8'h00;
		14'h39d6:	ff_dbi <= 8'h00;
		14'h39d7:	ff_dbi <= 8'h00;
		14'h39d8:	ff_dbi <= 8'h00;
		14'h39d9:	ff_dbi <= 8'h00;
		14'h39da:	ff_dbi <= 8'h00;
		14'h39db:	ff_dbi <= 8'h00;
		14'h39dc:	ff_dbi <= 8'h00;
		14'h39dd:	ff_dbi <= 8'h00;
		14'h39de:	ff_dbi <= 8'h00;
		14'h39df:	ff_dbi <= 8'h00;
		14'h39e0:	ff_dbi <= 8'h00;
		14'h39e1:	ff_dbi <= 8'h00;
		14'h39e2:	ff_dbi <= 8'h00;
		14'h39e3:	ff_dbi <= 8'h00;
		14'h39e4:	ff_dbi <= 8'h00;
		14'h39e5:	ff_dbi <= 8'h00;
		14'h39e6:	ff_dbi <= 8'h00;
		14'h39e7:	ff_dbi <= 8'h00;
		14'h39e8:	ff_dbi <= 8'h00;
		14'h39e9:	ff_dbi <= 8'h00;
		14'h39ea:	ff_dbi <= 8'h00;
		14'h39eb:	ff_dbi <= 8'h00;
		14'h39ec:	ff_dbi <= 8'h00;
		14'h39ed:	ff_dbi <= 8'h00;
		14'h39ee:	ff_dbi <= 8'h00;
		14'h39ef:	ff_dbi <= 8'h00;
		14'h39f0:	ff_dbi <= 8'h00;
		14'h39f1:	ff_dbi <= 8'h00;
		14'h39f2:	ff_dbi <= 8'h00;
		14'h39f3:	ff_dbi <= 8'h00;
		14'h39f4:	ff_dbi <= 8'h00;
		14'h39f5:	ff_dbi <= 8'h00;
		14'h39f6:	ff_dbi <= 8'h00;
		14'h39f7:	ff_dbi <= 8'h00;
		14'h39f8:	ff_dbi <= 8'h00;
		14'h39f9:	ff_dbi <= 8'h00;
		14'h39fa:	ff_dbi <= 8'h00;
		14'h39fb:	ff_dbi <= 8'h00;
		14'h39fc:	ff_dbi <= 8'h00;
		14'h39fd:	ff_dbi <= 8'h00;
		14'h39fe:	ff_dbi <= 8'h00;
		14'h39ff:	ff_dbi <= 8'h00;
		14'h3a00:	ff_dbi <= 8'h00;
		14'h3a01:	ff_dbi <= 8'h00;
		14'h3a02:	ff_dbi <= 8'h00;
		14'h3a03:	ff_dbi <= 8'h00;
		14'h3a04:	ff_dbi <= 8'h00;
		14'h3a05:	ff_dbi <= 8'h00;
		14'h3a06:	ff_dbi <= 8'h00;
		14'h3a07:	ff_dbi <= 8'h00;
		14'h3a08:	ff_dbi <= 8'h00;
		14'h3a09:	ff_dbi <= 8'h00;
		14'h3a0a:	ff_dbi <= 8'h00;
		14'h3a0b:	ff_dbi <= 8'h00;
		14'h3a0c:	ff_dbi <= 8'h00;
		14'h3a0d:	ff_dbi <= 8'h00;
		14'h3a0e:	ff_dbi <= 8'h00;
		14'h3a0f:	ff_dbi <= 8'h00;
		14'h3a10:	ff_dbi <= 8'h00;
		14'h3a11:	ff_dbi <= 8'h00;
		14'h3a12:	ff_dbi <= 8'h00;
		14'h3a13:	ff_dbi <= 8'h00;
		14'h3a14:	ff_dbi <= 8'h00;
		14'h3a15:	ff_dbi <= 8'h00;
		14'h3a16:	ff_dbi <= 8'h00;
		14'h3a17:	ff_dbi <= 8'h00;
		14'h3a18:	ff_dbi <= 8'h00;
		14'h3a19:	ff_dbi <= 8'h00;
		14'h3a1a:	ff_dbi <= 8'h00;
		14'h3a1b:	ff_dbi <= 8'h00;
		14'h3a1c:	ff_dbi <= 8'h00;
		14'h3a1d:	ff_dbi <= 8'h00;
		14'h3a1e:	ff_dbi <= 8'h00;
		14'h3a1f:	ff_dbi <= 8'h00;
		14'h3a20:	ff_dbi <= 8'h00;
		14'h3a21:	ff_dbi <= 8'h00;
		14'h3a22:	ff_dbi <= 8'h00;
		14'h3a23:	ff_dbi <= 8'h00;
		14'h3a24:	ff_dbi <= 8'h00;
		14'h3a25:	ff_dbi <= 8'h00;
		14'h3a26:	ff_dbi <= 8'h00;
		14'h3a27:	ff_dbi <= 8'h00;
		14'h3a28:	ff_dbi <= 8'h00;
		14'h3a29:	ff_dbi <= 8'h00;
		14'h3a2a:	ff_dbi <= 8'h00;
		14'h3a2b:	ff_dbi <= 8'h00;
		14'h3a2c:	ff_dbi <= 8'h00;
		14'h3a2d:	ff_dbi <= 8'h00;
		14'h3a2e:	ff_dbi <= 8'h00;
		14'h3a2f:	ff_dbi <= 8'h00;
		14'h3a30:	ff_dbi <= 8'h00;
		14'h3a31:	ff_dbi <= 8'h00;
		14'h3a32:	ff_dbi <= 8'h00;
		14'h3a33:	ff_dbi <= 8'h00;
		14'h3a34:	ff_dbi <= 8'h00;
		14'h3a35:	ff_dbi <= 8'h00;
		14'h3a36:	ff_dbi <= 8'h00;
		14'h3a37:	ff_dbi <= 8'h00;
		14'h3a38:	ff_dbi <= 8'h00;
		14'h3a39:	ff_dbi <= 8'h00;
		14'h3a3a:	ff_dbi <= 8'h00;
		14'h3a3b:	ff_dbi <= 8'h00;
		14'h3a3c:	ff_dbi <= 8'h00;
		14'h3a3d:	ff_dbi <= 8'h00;
		14'h3a3e:	ff_dbi <= 8'h00;
		14'h3a3f:	ff_dbi <= 8'h00;
		14'h3a40:	ff_dbi <= 8'h00;
		14'h3a41:	ff_dbi <= 8'h00;
		14'h3a42:	ff_dbi <= 8'h00;
		14'h3a43:	ff_dbi <= 8'h00;
		14'h3a44:	ff_dbi <= 8'h00;
		14'h3a45:	ff_dbi <= 8'h00;
		14'h3a46:	ff_dbi <= 8'h00;
		14'h3a47:	ff_dbi <= 8'h00;
		14'h3a48:	ff_dbi <= 8'h00;
		14'h3a49:	ff_dbi <= 8'h00;
		14'h3a4a:	ff_dbi <= 8'h00;
		14'h3a4b:	ff_dbi <= 8'h00;
		14'h3a4c:	ff_dbi <= 8'h00;
		14'h3a4d:	ff_dbi <= 8'h00;
		14'h3a4e:	ff_dbi <= 8'h00;
		14'h3a4f:	ff_dbi <= 8'h00;
		14'h3a50:	ff_dbi <= 8'h00;
		14'h3a51:	ff_dbi <= 8'h00;
		14'h3a52:	ff_dbi <= 8'h00;
		14'h3a53:	ff_dbi <= 8'h00;
		14'h3a54:	ff_dbi <= 8'h00;
		14'h3a55:	ff_dbi <= 8'h00;
		14'h3a56:	ff_dbi <= 8'h00;
		14'h3a57:	ff_dbi <= 8'h00;
		14'h3a58:	ff_dbi <= 8'h00;
		14'h3a59:	ff_dbi <= 8'h00;
		14'h3a5a:	ff_dbi <= 8'h00;
		14'h3a5b:	ff_dbi <= 8'h00;
		14'h3a5c:	ff_dbi <= 8'h00;
		14'h3a5d:	ff_dbi <= 8'h00;
		14'h3a5e:	ff_dbi <= 8'h00;
		14'h3a5f:	ff_dbi <= 8'h00;
		14'h3a60:	ff_dbi <= 8'h00;
		14'h3a61:	ff_dbi <= 8'h00;
		14'h3a62:	ff_dbi <= 8'h00;
		14'h3a63:	ff_dbi <= 8'h00;
		14'h3a64:	ff_dbi <= 8'h00;
		14'h3a65:	ff_dbi <= 8'h00;
		14'h3a66:	ff_dbi <= 8'h00;
		14'h3a67:	ff_dbi <= 8'h00;
		14'h3a68:	ff_dbi <= 8'h00;
		14'h3a69:	ff_dbi <= 8'h00;
		14'h3a6a:	ff_dbi <= 8'h00;
		14'h3a6b:	ff_dbi <= 8'h00;
		14'h3a6c:	ff_dbi <= 8'h00;
		14'h3a6d:	ff_dbi <= 8'h00;
		14'h3a6e:	ff_dbi <= 8'h00;
		14'h3a6f:	ff_dbi <= 8'h00;
		14'h3a70:	ff_dbi <= 8'h00;
		14'h3a71:	ff_dbi <= 8'h00;
		14'h3a72:	ff_dbi <= 8'h00;
		14'h3a73:	ff_dbi <= 8'h00;
		14'h3a74:	ff_dbi <= 8'h00;
		14'h3a75:	ff_dbi <= 8'h00;
		14'h3a76:	ff_dbi <= 8'h00;
		14'h3a77:	ff_dbi <= 8'h00;
		14'h3a78:	ff_dbi <= 8'h00;
		14'h3a79:	ff_dbi <= 8'h00;
		14'h3a7a:	ff_dbi <= 8'h00;
		14'h3a7b:	ff_dbi <= 8'h00;
		14'h3a7c:	ff_dbi <= 8'h00;
		14'h3a7d:	ff_dbi <= 8'h00;
		14'h3a7e:	ff_dbi <= 8'h00;
		14'h3a7f:	ff_dbi <= 8'h00;
		14'h3a80:	ff_dbi <= 8'h00;
		14'h3a81:	ff_dbi <= 8'h00;
		14'h3a82:	ff_dbi <= 8'h00;
		14'h3a83:	ff_dbi <= 8'h00;
		14'h3a84:	ff_dbi <= 8'h00;
		14'h3a85:	ff_dbi <= 8'h00;
		14'h3a86:	ff_dbi <= 8'h00;
		14'h3a87:	ff_dbi <= 8'h00;
		14'h3a88:	ff_dbi <= 8'h00;
		14'h3a89:	ff_dbi <= 8'h00;
		14'h3a8a:	ff_dbi <= 8'h00;
		14'h3a8b:	ff_dbi <= 8'h00;
		14'h3a8c:	ff_dbi <= 8'h00;
		14'h3a8d:	ff_dbi <= 8'h00;
		14'h3a8e:	ff_dbi <= 8'h00;
		14'h3a8f:	ff_dbi <= 8'h00;
		14'h3a90:	ff_dbi <= 8'h00;
		14'h3a91:	ff_dbi <= 8'h00;
		14'h3a92:	ff_dbi <= 8'h00;
		14'h3a93:	ff_dbi <= 8'h00;
		14'h3a94:	ff_dbi <= 8'h00;
		14'h3a95:	ff_dbi <= 8'h00;
		14'h3a96:	ff_dbi <= 8'h00;
		14'h3a97:	ff_dbi <= 8'h00;
		14'h3a98:	ff_dbi <= 8'h00;
		14'h3a99:	ff_dbi <= 8'h00;
		14'h3a9a:	ff_dbi <= 8'h00;
		14'h3a9b:	ff_dbi <= 8'h00;
		14'h3a9c:	ff_dbi <= 8'h00;
		14'h3a9d:	ff_dbi <= 8'h00;
		14'h3a9e:	ff_dbi <= 8'h00;
		14'h3a9f:	ff_dbi <= 8'h00;
		14'h3aa0:	ff_dbi <= 8'h00;
		14'h3aa1:	ff_dbi <= 8'h00;
		14'h3aa2:	ff_dbi <= 8'h00;
		14'h3aa3:	ff_dbi <= 8'h00;
		14'h3aa4:	ff_dbi <= 8'h00;
		14'h3aa5:	ff_dbi <= 8'h00;
		14'h3aa6:	ff_dbi <= 8'h00;
		14'h3aa7:	ff_dbi <= 8'h00;
		14'h3aa8:	ff_dbi <= 8'h00;
		14'h3aa9:	ff_dbi <= 8'h00;
		14'h3aaa:	ff_dbi <= 8'h00;
		14'h3aab:	ff_dbi <= 8'h00;
		14'h3aac:	ff_dbi <= 8'h00;
		14'h3aad:	ff_dbi <= 8'h00;
		14'h3aae:	ff_dbi <= 8'h00;
		14'h3aaf:	ff_dbi <= 8'h00;
		14'h3ab0:	ff_dbi <= 8'h00;
		14'h3ab1:	ff_dbi <= 8'h00;
		14'h3ab2:	ff_dbi <= 8'h00;
		14'h3ab3:	ff_dbi <= 8'h00;
		14'h3ab4:	ff_dbi <= 8'h00;
		14'h3ab5:	ff_dbi <= 8'h00;
		14'h3ab6:	ff_dbi <= 8'h00;
		14'h3ab7:	ff_dbi <= 8'h00;
		14'h3ab8:	ff_dbi <= 8'h00;
		14'h3ab9:	ff_dbi <= 8'h00;
		14'h3aba:	ff_dbi <= 8'h00;
		14'h3abb:	ff_dbi <= 8'h00;
		14'h3abc:	ff_dbi <= 8'h00;
		14'h3abd:	ff_dbi <= 8'h00;
		14'h3abe:	ff_dbi <= 8'h00;
		14'h3abf:	ff_dbi <= 8'h00;
		14'h3ac0:	ff_dbi <= 8'h00;
		14'h3ac1:	ff_dbi <= 8'h00;
		14'h3ac2:	ff_dbi <= 8'h00;
		14'h3ac3:	ff_dbi <= 8'h00;
		14'h3ac4:	ff_dbi <= 8'h00;
		14'h3ac5:	ff_dbi <= 8'h00;
		14'h3ac6:	ff_dbi <= 8'h00;
		14'h3ac7:	ff_dbi <= 8'h00;
		14'h3ac8:	ff_dbi <= 8'h00;
		14'h3ac9:	ff_dbi <= 8'h00;
		14'h3aca:	ff_dbi <= 8'h00;
		14'h3acb:	ff_dbi <= 8'h00;
		14'h3acc:	ff_dbi <= 8'h00;
		14'h3acd:	ff_dbi <= 8'h00;
		14'h3ace:	ff_dbi <= 8'h00;
		14'h3acf:	ff_dbi <= 8'h00;
		14'h3ad0:	ff_dbi <= 8'h00;
		14'h3ad1:	ff_dbi <= 8'h00;
		14'h3ad2:	ff_dbi <= 8'h00;
		14'h3ad3:	ff_dbi <= 8'h00;
		14'h3ad4:	ff_dbi <= 8'h00;
		14'h3ad5:	ff_dbi <= 8'h00;
		14'h3ad6:	ff_dbi <= 8'h00;
		14'h3ad7:	ff_dbi <= 8'h00;
		14'h3ad8:	ff_dbi <= 8'h00;
		14'h3ad9:	ff_dbi <= 8'h00;
		14'h3ada:	ff_dbi <= 8'h00;
		14'h3adb:	ff_dbi <= 8'h00;
		14'h3adc:	ff_dbi <= 8'h00;
		14'h3add:	ff_dbi <= 8'h00;
		14'h3ade:	ff_dbi <= 8'h00;
		14'h3adf:	ff_dbi <= 8'h00;
		14'h3ae0:	ff_dbi <= 8'h00;
		14'h3ae1:	ff_dbi <= 8'h00;
		14'h3ae2:	ff_dbi <= 8'h00;
		14'h3ae3:	ff_dbi <= 8'h00;
		14'h3ae4:	ff_dbi <= 8'h00;
		14'h3ae5:	ff_dbi <= 8'h00;
		14'h3ae6:	ff_dbi <= 8'h00;
		14'h3ae7:	ff_dbi <= 8'h00;
		14'h3ae8:	ff_dbi <= 8'h00;
		14'h3ae9:	ff_dbi <= 8'h00;
		14'h3aea:	ff_dbi <= 8'h00;
		14'h3aeb:	ff_dbi <= 8'h00;
		14'h3aec:	ff_dbi <= 8'h00;
		14'h3aed:	ff_dbi <= 8'h00;
		14'h3aee:	ff_dbi <= 8'h00;
		14'h3aef:	ff_dbi <= 8'h00;
		14'h3af0:	ff_dbi <= 8'h00;
		14'h3af1:	ff_dbi <= 8'h00;
		14'h3af2:	ff_dbi <= 8'h00;
		14'h3af3:	ff_dbi <= 8'h00;
		14'h3af4:	ff_dbi <= 8'h00;
		14'h3af5:	ff_dbi <= 8'h00;
		14'h3af6:	ff_dbi <= 8'h00;
		14'h3af7:	ff_dbi <= 8'h00;
		14'h3af8:	ff_dbi <= 8'h00;
		14'h3af9:	ff_dbi <= 8'h00;
		14'h3afa:	ff_dbi <= 8'h00;
		14'h3afb:	ff_dbi <= 8'h00;
		14'h3afc:	ff_dbi <= 8'h00;
		14'h3afd:	ff_dbi <= 8'h00;
		14'h3afe:	ff_dbi <= 8'h00;
		14'h3aff:	ff_dbi <= 8'h00;
		14'h3b00:	ff_dbi <= 8'h00;
		14'h3b01:	ff_dbi <= 8'h00;
		14'h3b02:	ff_dbi <= 8'h00;
		14'h3b03:	ff_dbi <= 8'h00;
		14'h3b04:	ff_dbi <= 8'h00;
		14'h3b05:	ff_dbi <= 8'h00;
		14'h3b06:	ff_dbi <= 8'h00;
		14'h3b07:	ff_dbi <= 8'h00;
		14'h3b08:	ff_dbi <= 8'h00;
		14'h3b09:	ff_dbi <= 8'h00;
		14'h3b0a:	ff_dbi <= 8'h00;
		14'h3b0b:	ff_dbi <= 8'h00;
		14'h3b0c:	ff_dbi <= 8'h00;
		14'h3b0d:	ff_dbi <= 8'h00;
		14'h3b0e:	ff_dbi <= 8'h00;
		14'h3b0f:	ff_dbi <= 8'h00;
		14'h3b10:	ff_dbi <= 8'h00;
		14'h3b11:	ff_dbi <= 8'h00;
		14'h3b12:	ff_dbi <= 8'h00;
		14'h3b13:	ff_dbi <= 8'h00;
		14'h3b14:	ff_dbi <= 8'h00;
		14'h3b15:	ff_dbi <= 8'h00;
		14'h3b16:	ff_dbi <= 8'h00;
		14'h3b17:	ff_dbi <= 8'h00;
		14'h3b18:	ff_dbi <= 8'h00;
		14'h3b19:	ff_dbi <= 8'h00;
		14'h3b1a:	ff_dbi <= 8'h00;
		14'h3b1b:	ff_dbi <= 8'h00;
		14'h3b1c:	ff_dbi <= 8'h00;
		14'h3b1d:	ff_dbi <= 8'h00;
		14'h3b1e:	ff_dbi <= 8'h00;
		14'h3b1f:	ff_dbi <= 8'h00;
		14'h3b20:	ff_dbi <= 8'h00;
		14'h3b21:	ff_dbi <= 8'h00;
		14'h3b22:	ff_dbi <= 8'h00;
		14'h3b23:	ff_dbi <= 8'h00;
		14'h3b24:	ff_dbi <= 8'h00;
		14'h3b25:	ff_dbi <= 8'h00;
		14'h3b26:	ff_dbi <= 8'h00;
		14'h3b27:	ff_dbi <= 8'h00;
		14'h3b28:	ff_dbi <= 8'h00;
		14'h3b29:	ff_dbi <= 8'h00;
		14'h3b2a:	ff_dbi <= 8'h00;
		14'h3b2b:	ff_dbi <= 8'h00;
		14'h3b2c:	ff_dbi <= 8'h00;
		14'h3b2d:	ff_dbi <= 8'h00;
		14'h3b2e:	ff_dbi <= 8'h00;
		14'h3b2f:	ff_dbi <= 8'h00;
		14'h3b30:	ff_dbi <= 8'h00;
		14'h3b31:	ff_dbi <= 8'h00;
		14'h3b32:	ff_dbi <= 8'h00;
		14'h3b33:	ff_dbi <= 8'h00;
		14'h3b34:	ff_dbi <= 8'h00;
		14'h3b35:	ff_dbi <= 8'h00;
		14'h3b36:	ff_dbi <= 8'h00;
		14'h3b37:	ff_dbi <= 8'h00;
		14'h3b38:	ff_dbi <= 8'h00;
		14'h3b39:	ff_dbi <= 8'h00;
		14'h3b3a:	ff_dbi <= 8'h00;
		14'h3b3b:	ff_dbi <= 8'h00;
		14'h3b3c:	ff_dbi <= 8'h00;
		14'h3b3d:	ff_dbi <= 8'h00;
		14'h3b3e:	ff_dbi <= 8'h00;
		14'h3b3f:	ff_dbi <= 8'h00;
		14'h3b40:	ff_dbi <= 8'h00;
		14'h3b41:	ff_dbi <= 8'h00;
		14'h3b42:	ff_dbi <= 8'h00;
		14'h3b43:	ff_dbi <= 8'h00;
		14'h3b44:	ff_dbi <= 8'h00;
		14'h3b45:	ff_dbi <= 8'h00;
		14'h3b46:	ff_dbi <= 8'h00;
		14'h3b47:	ff_dbi <= 8'h00;
		14'h3b48:	ff_dbi <= 8'h00;
		14'h3b49:	ff_dbi <= 8'h00;
		14'h3b4a:	ff_dbi <= 8'h00;
		14'h3b4b:	ff_dbi <= 8'h00;
		14'h3b4c:	ff_dbi <= 8'h00;
		14'h3b4d:	ff_dbi <= 8'h00;
		14'h3b4e:	ff_dbi <= 8'h00;
		14'h3b4f:	ff_dbi <= 8'h00;
		14'h3b50:	ff_dbi <= 8'h00;
		14'h3b51:	ff_dbi <= 8'h00;
		14'h3b52:	ff_dbi <= 8'h00;
		14'h3b53:	ff_dbi <= 8'h00;
		14'h3b54:	ff_dbi <= 8'h00;
		14'h3b55:	ff_dbi <= 8'h00;
		14'h3b56:	ff_dbi <= 8'h00;
		14'h3b57:	ff_dbi <= 8'h00;
		14'h3b58:	ff_dbi <= 8'h00;
		14'h3b59:	ff_dbi <= 8'h00;
		14'h3b5a:	ff_dbi <= 8'h00;
		14'h3b5b:	ff_dbi <= 8'h00;
		14'h3b5c:	ff_dbi <= 8'h00;
		14'h3b5d:	ff_dbi <= 8'h00;
		14'h3b5e:	ff_dbi <= 8'h00;
		14'h3b5f:	ff_dbi <= 8'h00;
		14'h3b60:	ff_dbi <= 8'h00;
		14'h3b61:	ff_dbi <= 8'h00;
		14'h3b62:	ff_dbi <= 8'h00;
		14'h3b63:	ff_dbi <= 8'h00;
		14'h3b64:	ff_dbi <= 8'h00;
		14'h3b65:	ff_dbi <= 8'h00;
		14'h3b66:	ff_dbi <= 8'h00;
		14'h3b67:	ff_dbi <= 8'h00;
		14'h3b68:	ff_dbi <= 8'h00;
		14'h3b69:	ff_dbi <= 8'h00;
		14'h3b6a:	ff_dbi <= 8'h00;
		14'h3b6b:	ff_dbi <= 8'h00;
		14'h3b6c:	ff_dbi <= 8'h00;
		14'h3b6d:	ff_dbi <= 8'h00;
		14'h3b6e:	ff_dbi <= 8'h00;
		14'h3b6f:	ff_dbi <= 8'h00;
		14'h3b70:	ff_dbi <= 8'h00;
		14'h3b71:	ff_dbi <= 8'h00;
		14'h3b72:	ff_dbi <= 8'h00;
		14'h3b73:	ff_dbi <= 8'h00;
		14'h3b74:	ff_dbi <= 8'h00;
		14'h3b75:	ff_dbi <= 8'h00;
		14'h3b76:	ff_dbi <= 8'h00;
		14'h3b77:	ff_dbi <= 8'h00;
		14'h3b78:	ff_dbi <= 8'h00;
		14'h3b79:	ff_dbi <= 8'h00;
		14'h3b7a:	ff_dbi <= 8'h00;
		14'h3b7b:	ff_dbi <= 8'h00;
		14'h3b7c:	ff_dbi <= 8'h00;
		14'h3b7d:	ff_dbi <= 8'h00;
		14'h3b7e:	ff_dbi <= 8'h00;
		14'h3b7f:	ff_dbi <= 8'h00;
		14'h3b80:	ff_dbi <= 8'h00;
		14'h3b81:	ff_dbi <= 8'h00;
		14'h3b82:	ff_dbi <= 8'h00;
		14'h3b83:	ff_dbi <= 8'h00;
		14'h3b84:	ff_dbi <= 8'h00;
		14'h3b85:	ff_dbi <= 8'h00;
		14'h3b86:	ff_dbi <= 8'h00;
		14'h3b87:	ff_dbi <= 8'h00;
		14'h3b88:	ff_dbi <= 8'h00;
		14'h3b89:	ff_dbi <= 8'h00;
		14'h3b8a:	ff_dbi <= 8'h00;
		14'h3b8b:	ff_dbi <= 8'h00;
		14'h3b8c:	ff_dbi <= 8'h00;
		14'h3b8d:	ff_dbi <= 8'h00;
		14'h3b8e:	ff_dbi <= 8'h00;
		14'h3b8f:	ff_dbi <= 8'h00;
		14'h3b90:	ff_dbi <= 8'h00;
		14'h3b91:	ff_dbi <= 8'h00;
		14'h3b92:	ff_dbi <= 8'h00;
		14'h3b93:	ff_dbi <= 8'h00;
		14'h3b94:	ff_dbi <= 8'h00;
		14'h3b95:	ff_dbi <= 8'h00;
		14'h3b96:	ff_dbi <= 8'h00;
		14'h3b97:	ff_dbi <= 8'h00;
		14'h3b98:	ff_dbi <= 8'h00;
		14'h3b99:	ff_dbi <= 8'h00;
		14'h3b9a:	ff_dbi <= 8'h00;
		14'h3b9b:	ff_dbi <= 8'h00;
		14'h3b9c:	ff_dbi <= 8'h00;
		14'h3b9d:	ff_dbi <= 8'h00;
		14'h3b9e:	ff_dbi <= 8'h00;
		14'h3b9f:	ff_dbi <= 8'h00;
		14'h3ba0:	ff_dbi <= 8'h00;
		14'h3ba1:	ff_dbi <= 8'h00;
		14'h3ba2:	ff_dbi <= 8'h00;
		14'h3ba3:	ff_dbi <= 8'h00;
		14'h3ba4:	ff_dbi <= 8'h00;
		14'h3ba5:	ff_dbi <= 8'h00;
		14'h3ba6:	ff_dbi <= 8'h00;
		14'h3ba7:	ff_dbi <= 8'h00;
		14'h3ba8:	ff_dbi <= 8'h00;
		14'h3ba9:	ff_dbi <= 8'h00;
		14'h3baa:	ff_dbi <= 8'h00;
		14'h3bab:	ff_dbi <= 8'h00;
		14'h3bac:	ff_dbi <= 8'h00;
		14'h3bad:	ff_dbi <= 8'h00;
		14'h3bae:	ff_dbi <= 8'h00;
		14'h3baf:	ff_dbi <= 8'h00;
		14'h3bb0:	ff_dbi <= 8'h00;
		14'h3bb1:	ff_dbi <= 8'h00;
		14'h3bb2:	ff_dbi <= 8'h00;
		14'h3bb3:	ff_dbi <= 8'h00;
		14'h3bb4:	ff_dbi <= 8'h00;
		14'h3bb5:	ff_dbi <= 8'h00;
		14'h3bb6:	ff_dbi <= 8'h00;
		14'h3bb7:	ff_dbi <= 8'h00;
		14'h3bb8:	ff_dbi <= 8'h00;
		14'h3bb9:	ff_dbi <= 8'h00;
		14'h3bba:	ff_dbi <= 8'h00;
		14'h3bbb:	ff_dbi <= 8'h00;
		14'h3bbc:	ff_dbi <= 8'h00;
		14'h3bbd:	ff_dbi <= 8'h00;
		14'h3bbe:	ff_dbi <= 8'h00;
		14'h3bbf:	ff_dbi <= 8'h00;
		14'h3bc0:	ff_dbi <= 8'h00;
		14'h3bc1:	ff_dbi <= 8'h00;
		14'h3bc2:	ff_dbi <= 8'h00;
		14'h3bc3:	ff_dbi <= 8'h00;
		14'h3bc4:	ff_dbi <= 8'h00;
		14'h3bc5:	ff_dbi <= 8'h00;
		14'h3bc6:	ff_dbi <= 8'h00;
		14'h3bc7:	ff_dbi <= 8'h00;
		14'h3bc8:	ff_dbi <= 8'h00;
		14'h3bc9:	ff_dbi <= 8'h00;
		14'h3bca:	ff_dbi <= 8'h00;
		14'h3bcb:	ff_dbi <= 8'h00;
		14'h3bcc:	ff_dbi <= 8'h00;
		14'h3bcd:	ff_dbi <= 8'h00;
		14'h3bce:	ff_dbi <= 8'h00;
		14'h3bcf:	ff_dbi <= 8'h00;
		14'h3bd0:	ff_dbi <= 8'h00;
		14'h3bd1:	ff_dbi <= 8'h00;
		14'h3bd2:	ff_dbi <= 8'h00;
		14'h3bd3:	ff_dbi <= 8'h00;
		14'h3bd4:	ff_dbi <= 8'h00;
		14'h3bd5:	ff_dbi <= 8'h00;
		14'h3bd6:	ff_dbi <= 8'h00;
		14'h3bd7:	ff_dbi <= 8'h00;
		14'h3bd8:	ff_dbi <= 8'h00;
		14'h3bd9:	ff_dbi <= 8'h00;
		14'h3bda:	ff_dbi <= 8'h00;
		14'h3bdb:	ff_dbi <= 8'h00;
		14'h3bdc:	ff_dbi <= 8'h00;
		14'h3bdd:	ff_dbi <= 8'h00;
		14'h3bde:	ff_dbi <= 8'h00;
		14'h3bdf:	ff_dbi <= 8'h00;
		14'h3be0:	ff_dbi <= 8'h00;
		14'h3be1:	ff_dbi <= 8'h00;
		14'h3be2:	ff_dbi <= 8'h00;
		14'h3be3:	ff_dbi <= 8'h00;
		14'h3be4:	ff_dbi <= 8'h00;
		14'h3be5:	ff_dbi <= 8'h00;
		14'h3be6:	ff_dbi <= 8'h00;
		14'h3be7:	ff_dbi <= 8'h00;
		14'h3be8:	ff_dbi <= 8'h00;
		14'h3be9:	ff_dbi <= 8'h00;
		14'h3bea:	ff_dbi <= 8'h00;
		14'h3beb:	ff_dbi <= 8'h00;
		14'h3bec:	ff_dbi <= 8'h00;
		14'h3bed:	ff_dbi <= 8'h00;
		14'h3bee:	ff_dbi <= 8'h00;
		14'h3bef:	ff_dbi <= 8'h00;
		14'h3bf0:	ff_dbi <= 8'h00;
		14'h3bf1:	ff_dbi <= 8'h00;
		14'h3bf2:	ff_dbi <= 8'h00;
		14'h3bf3:	ff_dbi <= 8'h00;
		14'h3bf4:	ff_dbi <= 8'h00;
		14'h3bf5:	ff_dbi <= 8'h00;
		14'h3bf6:	ff_dbi <= 8'h00;
		14'h3bf7:	ff_dbi <= 8'h00;
		14'h3bf8:	ff_dbi <= 8'h00;
		14'h3bf9:	ff_dbi <= 8'h00;
		14'h3bfa:	ff_dbi <= 8'h00;
		14'h3bfb:	ff_dbi <= 8'h00;
		14'h3bfc:	ff_dbi <= 8'h00;
		14'h3bfd:	ff_dbi <= 8'h00;
		14'h3bfe:	ff_dbi <= 8'h00;
		14'h3bff:	ff_dbi <= 8'h00;
		14'h3c00:	ff_dbi <= 8'h00;
		14'h3c01:	ff_dbi <= 8'h00;
		14'h3c02:	ff_dbi <= 8'h00;
		14'h3c03:	ff_dbi <= 8'h00;
		14'h3c04:	ff_dbi <= 8'h00;
		14'h3c05:	ff_dbi <= 8'h00;
		14'h3c06:	ff_dbi <= 8'h00;
		14'h3c07:	ff_dbi <= 8'h00;
		14'h3c08:	ff_dbi <= 8'h00;
		14'h3c09:	ff_dbi <= 8'h00;
		14'h3c0a:	ff_dbi <= 8'h00;
		14'h3c0b:	ff_dbi <= 8'h00;
		14'h3c0c:	ff_dbi <= 8'h00;
		14'h3c0d:	ff_dbi <= 8'h00;
		14'h3c0e:	ff_dbi <= 8'h00;
		14'h3c0f:	ff_dbi <= 8'h00;
		14'h3c10:	ff_dbi <= 8'h00;
		14'h3c11:	ff_dbi <= 8'h00;
		14'h3c12:	ff_dbi <= 8'h00;
		14'h3c13:	ff_dbi <= 8'h00;
		14'h3c14:	ff_dbi <= 8'h00;
		14'h3c15:	ff_dbi <= 8'h00;
		14'h3c16:	ff_dbi <= 8'h00;
		14'h3c17:	ff_dbi <= 8'h00;
		14'h3c18:	ff_dbi <= 8'h00;
		14'h3c19:	ff_dbi <= 8'h00;
		14'h3c1a:	ff_dbi <= 8'h00;
		14'h3c1b:	ff_dbi <= 8'h00;
		14'h3c1c:	ff_dbi <= 8'h00;
		14'h3c1d:	ff_dbi <= 8'h00;
		14'h3c1e:	ff_dbi <= 8'h00;
		14'h3c1f:	ff_dbi <= 8'h00;
		14'h3c20:	ff_dbi <= 8'h00;
		14'h3c21:	ff_dbi <= 8'h00;
		14'h3c22:	ff_dbi <= 8'h00;
		14'h3c23:	ff_dbi <= 8'h00;
		14'h3c24:	ff_dbi <= 8'h00;
		14'h3c25:	ff_dbi <= 8'h00;
		14'h3c26:	ff_dbi <= 8'h00;
		14'h3c27:	ff_dbi <= 8'h00;
		14'h3c28:	ff_dbi <= 8'h00;
		14'h3c29:	ff_dbi <= 8'h00;
		14'h3c2a:	ff_dbi <= 8'h00;
		14'h3c2b:	ff_dbi <= 8'h00;
		14'h3c2c:	ff_dbi <= 8'h00;
		14'h3c2d:	ff_dbi <= 8'h00;
		14'h3c2e:	ff_dbi <= 8'h00;
		14'h3c2f:	ff_dbi <= 8'h00;
		14'h3c30:	ff_dbi <= 8'h00;
		14'h3c31:	ff_dbi <= 8'h00;
		14'h3c32:	ff_dbi <= 8'h00;
		14'h3c33:	ff_dbi <= 8'h00;
		14'h3c34:	ff_dbi <= 8'h00;
		14'h3c35:	ff_dbi <= 8'h00;
		14'h3c36:	ff_dbi <= 8'h00;
		14'h3c37:	ff_dbi <= 8'h00;
		14'h3c38:	ff_dbi <= 8'h00;
		14'h3c39:	ff_dbi <= 8'h00;
		14'h3c3a:	ff_dbi <= 8'h00;
		14'h3c3b:	ff_dbi <= 8'h00;
		14'h3c3c:	ff_dbi <= 8'h00;
		14'h3c3d:	ff_dbi <= 8'h00;
		14'h3c3e:	ff_dbi <= 8'h00;
		14'h3c3f:	ff_dbi <= 8'h00;
		14'h3c40:	ff_dbi <= 8'h00;
		14'h3c41:	ff_dbi <= 8'h00;
		14'h3c42:	ff_dbi <= 8'h00;
		14'h3c43:	ff_dbi <= 8'h00;
		14'h3c44:	ff_dbi <= 8'h00;
		14'h3c45:	ff_dbi <= 8'h00;
		14'h3c46:	ff_dbi <= 8'h00;
		14'h3c47:	ff_dbi <= 8'h00;
		14'h3c48:	ff_dbi <= 8'h00;
		14'h3c49:	ff_dbi <= 8'h00;
		14'h3c4a:	ff_dbi <= 8'h00;
		14'h3c4b:	ff_dbi <= 8'h00;
		14'h3c4c:	ff_dbi <= 8'h00;
		14'h3c4d:	ff_dbi <= 8'h00;
		14'h3c4e:	ff_dbi <= 8'h00;
		14'h3c4f:	ff_dbi <= 8'h00;
		14'h3c50:	ff_dbi <= 8'h00;
		14'h3c51:	ff_dbi <= 8'h00;
		14'h3c52:	ff_dbi <= 8'h00;
		14'h3c53:	ff_dbi <= 8'h00;
		14'h3c54:	ff_dbi <= 8'h00;
		14'h3c55:	ff_dbi <= 8'h00;
		14'h3c56:	ff_dbi <= 8'h00;
		14'h3c57:	ff_dbi <= 8'h00;
		14'h3c58:	ff_dbi <= 8'h00;
		14'h3c59:	ff_dbi <= 8'h00;
		14'h3c5a:	ff_dbi <= 8'h00;
		14'h3c5b:	ff_dbi <= 8'h00;
		14'h3c5c:	ff_dbi <= 8'h00;
		14'h3c5d:	ff_dbi <= 8'h00;
		14'h3c5e:	ff_dbi <= 8'h00;
		14'h3c5f:	ff_dbi <= 8'h00;
		14'h3c60:	ff_dbi <= 8'h00;
		14'h3c61:	ff_dbi <= 8'h00;
		14'h3c62:	ff_dbi <= 8'h00;
		14'h3c63:	ff_dbi <= 8'h00;
		14'h3c64:	ff_dbi <= 8'h00;
		14'h3c65:	ff_dbi <= 8'h00;
		14'h3c66:	ff_dbi <= 8'h00;
		14'h3c67:	ff_dbi <= 8'h00;
		14'h3c68:	ff_dbi <= 8'h00;
		14'h3c69:	ff_dbi <= 8'h00;
		14'h3c6a:	ff_dbi <= 8'h00;
		14'h3c6b:	ff_dbi <= 8'h00;
		14'h3c6c:	ff_dbi <= 8'h00;
		14'h3c6d:	ff_dbi <= 8'h00;
		14'h3c6e:	ff_dbi <= 8'h00;
		14'h3c6f:	ff_dbi <= 8'h00;
		14'h3c70:	ff_dbi <= 8'h00;
		14'h3c71:	ff_dbi <= 8'h00;
		14'h3c72:	ff_dbi <= 8'h00;
		14'h3c73:	ff_dbi <= 8'h00;
		14'h3c74:	ff_dbi <= 8'h00;
		14'h3c75:	ff_dbi <= 8'h00;
		14'h3c76:	ff_dbi <= 8'h00;
		14'h3c77:	ff_dbi <= 8'h00;
		14'h3c78:	ff_dbi <= 8'h00;
		14'h3c79:	ff_dbi <= 8'h00;
		14'h3c7a:	ff_dbi <= 8'h00;
		14'h3c7b:	ff_dbi <= 8'h00;
		14'h3c7c:	ff_dbi <= 8'h00;
		14'h3c7d:	ff_dbi <= 8'h00;
		14'h3c7e:	ff_dbi <= 8'h00;
		14'h3c7f:	ff_dbi <= 8'h00;
		14'h3c80:	ff_dbi <= 8'h00;
		14'h3c81:	ff_dbi <= 8'h00;
		14'h3c82:	ff_dbi <= 8'h00;
		14'h3c83:	ff_dbi <= 8'h00;
		14'h3c84:	ff_dbi <= 8'h00;
		14'h3c85:	ff_dbi <= 8'h00;
		14'h3c86:	ff_dbi <= 8'h00;
		14'h3c87:	ff_dbi <= 8'h00;
		14'h3c88:	ff_dbi <= 8'h00;
		14'h3c89:	ff_dbi <= 8'h00;
		14'h3c8a:	ff_dbi <= 8'h00;
		14'h3c8b:	ff_dbi <= 8'h00;
		14'h3c8c:	ff_dbi <= 8'h00;
		14'h3c8d:	ff_dbi <= 8'h00;
		14'h3c8e:	ff_dbi <= 8'h00;
		14'h3c8f:	ff_dbi <= 8'h00;
		14'h3c90:	ff_dbi <= 8'h00;
		14'h3c91:	ff_dbi <= 8'h00;
		14'h3c92:	ff_dbi <= 8'h00;
		14'h3c93:	ff_dbi <= 8'h00;
		14'h3c94:	ff_dbi <= 8'h00;
		14'h3c95:	ff_dbi <= 8'h00;
		14'h3c96:	ff_dbi <= 8'h00;
		14'h3c97:	ff_dbi <= 8'h00;
		14'h3c98:	ff_dbi <= 8'h00;
		14'h3c99:	ff_dbi <= 8'h00;
		14'h3c9a:	ff_dbi <= 8'h00;
		14'h3c9b:	ff_dbi <= 8'h00;
		14'h3c9c:	ff_dbi <= 8'h00;
		14'h3c9d:	ff_dbi <= 8'h00;
		14'h3c9e:	ff_dbi <= 8'h00;
		14'h3c9f:	ff_dbi <= 8'h00;
		14'h3ca0:	ff_dbi <= 8'h00;
		14'h3ca1:	ff_dbi <= 8'h00;
		14'h3ca2:	ff_dbi <= 8'h00;
		14'h3ca3:	ff_dbi <= 8'h00;
		14'h3ca4:	ff_dbi <= 8'h00;
		14'h3ca5:	ff_dbi <= 8'h00;
		14'h3ca6:	ff_dbi <= 8'h00;
		14'h3ca7:	ff_dbi <= 8'h00;
		14'h3ca8:	ff_dbi <= 8'h00;
		14'h3ca9:	ff_dbi <= 8'h00;
		14'h3caa:	ff_dbi <= 8'h00;
		14'h3cab:	ff_dbi <= 8'h00;
		14'h3cac:	ff_dbi <= 8'h00;
		14'h3cad:	ff_dbi <= 8'h00;
		14'h3cae:	ff_dbi <= 8'h00;
		14'h3caf:	ff_dbi <= 8'h00;
		14'h3cb0:	ff_dbi <= 8'h00;
		14'h3cb1:	ff_dbi <= 8'h00;
		14'h3cb2:	ff_dbi <= 8'h00;
		14'h3cb3:	ff_dbi <= 8'h00;
		14'h3cb4:	ff_dbi <= 8'h00;
		14'h3cb5:	ff_dbi <= 8'h00;
		14'h3cb6:	ff_dbi <= 8'h00;
		14'h3cb7:	ff_dbi <= 8'h00;
		14'h3cb8:	ff_dbi <= 8'h00;
		14'h3cb9:	ff_dbi <= 8'h00;
		14'h3cba:	ff_dbi <= 8'h00;
		14'h3cbb:	ff_dbi <= 8'h00;
		14'h3cbc:	ff_dbi <= 8'h00;
		14'h3cbd:	ff_dbi <= 8'h00;
		14'h3cbe:	ff_dbi <= 8'h00;
		14'h3cbf:	ff_dbi <= 8'h00;
		14'h3cc0:	ff_dbi <= 8'h00;
		14'h3cc1:	ff_dbi <= 8'h00;
		14'h3cc2:	ff_dbi <= 8'h00;
		14'h3cc3:	ff_dbi <= 8'h00;
		14'h3cc4:	ff_dbi <= 8'h00;
		14'h3cc5:	ff_dbi <= 8'h00;
		14'h3cc6:	ff_dbi <= 8'h00;
		14'h3cc7:	ff_dbi <= 8'h00;
		14'h3cc8:	ff_dbi <= 8'h00;
		14'h3cc9:	ff_dbi <= 8'h00;
		14'h3cca:	ff_dbi <= 8'h00;
		14'h3ccb:	ff_dbi <= 8'h00;
		14'h3ccc:	ff_dbi <= 8'h00;
		14'h3ccd:	ff_dbi <= 8'h00;
		14'h3cce:	ff_dbi <= 8'h00;
		14'h3ccf:	ff_dbi <= 8'h00;
		14'h3cd0:	ff_dbi <= 8'h00;
		14'h3cd1:	ff_dbi <= 8'h00;
		14'h3cd2:	ff_dbi <= 8'h00;
		14'h3cd3:	ff_dbi <= 8'h00;
		14'h3cd4:	ff_dbi <= 8'h00;
		14'h3cd5:	ff_dbi <= 8'h00;
		14'h3cd6:	ff_dbi <= 8'h00;
		14'h3cd7:	ff_dbi <= 8'h00;
		14'h3cd8:	ff_dbi <= 8'h00;
		14'h3cd9:	ff_dbi <= 8'h00;
		14'h3cda:	ff_dbi <= 8'h00;
		14'h3cdb:	ff_dbi <= 8'h00;
		14'h3cdc:	ff_dbi <= 8'h00;
		14'h3cdd:	ff_dbi <= 8'h00;
		14'h3cde:	ff_dbi <= 8'h00;
		14'h3cdf:	ff_dbi <= 8'h00;
		14'h3ce0:	ff_dbi <= 8'h00;
		14'h3ce1:	ff_dbi <= 8'h00;
		14'h3ce2:	ff_dbi <= 8'h00;
		14'h3ce3:	ff_dbi <= 8'h00;
		14'h3ce4:	ff_dbi <= 8'h00;
		14'h3ce5:	ff_dbi <= 8'h00;
		14'h3ce6:	ff_dbi <= 8'h00;
		14'h3ce7:	ff_dbi <= 8'h00;
		14'h3ce8:	ff_dbi <= 8'h00;
		14'h3ce9:	ff_dbi <= 8'h00;
		14'h3cea:	ff_dbi <= 8'h00;
		14'h3ceb:	ff_dbi <= 8'h00;
		14'h3cec:	ff_dbi <= 8'h00;
		14'h3ced:	ff_dbi <= 8'h00;
		14'h3cee:	ff_dbi <= 8'h00;
		14'h3cef:	ff_dbi <= 8'h00;
		14'h3cf0:	ff_dbi <= 8'h00;
		14'h3cf1:	ff_dbi <= 8'h00;
		14'h3cf2:	ff_dbi <= 8'h00;
		14'h3cf3:	ff_dbi <= 8'h00;
		14'h3cf4:	ff_dbi <= 8'h00;
		14'h3cf5:	ff_dbi <= 8'h00;
		14'h3cf6:	ff_dbi <= 8'h00;
		14'h3cf7:	ff_dbi <= 8'h00;
		14'h3cf8:	ff_dbi <= 8'h00;
		14'h3cf9:	ff_dbi <= 8'h00;
		14'h3cfa:	ff_dbi <= 8'h00;
		14'h3cfb:	ff_dbi <= 8'h00;
		14'h3cfc:	ff_dbi <= 8'h00;
		14'h3cfd:	ff_dbi <= 8'h00;
		14'h3cfe:	ff_dbi <= 8'h00;
		14'h3cff:	ff_dbi <= 8'h00;
		14'h3d00:	ff_dbi <= 8'h00;
		14'h3d01:	ff_dbi <= 8'h00;
		14'h3d02:	ff_dbi <= 8'h00;
		14'h3d03:	ff_dbi <= 8'h00;
		14'h3d04:	ff_dbi <= 8'h00;
		14'h3d05:	ff_dbi <= 8'h00;
		14'h3d06:	ff_dbi <= 8'h00;
		14'h3d07:	ff_dbi <= 8'h00;
		14'h3d08:	ff_dbi <= 8'h00;
		14'h3d09:	ff_dbi <= 8'h00;
		14'h3d0a:	ff_dbi <= 8'h00;
		14'h3d0b:	ff_dbi <= 8'h00;
		14'h3d0c:	ff_dbi <= 8'h00;
		14'h3d0d:	ff_dbi <= 8'h00;
		14'h3d0e:	ff_dbi <= 8'h00;
		14'h3d0f:	ff_dbi <= 8'h00;
		14'h3d10:	ff_dbi <= 8'h00;
		14'h3d11:	ff_dbi <= 8'h00;
		14'h3d12:	ff_dbi <= 8'h00;
		14'h3d13:	ff_dbi <= 8'h00;
		14'h3d14:	ff_dbi <= 8'h00;
		14'h3d15:	ff_dbi <= 8'h00;
		14'h3d16:	ff_dbi <= 8'h00;
		14'h3d17:	ff_dbi <= 8'h00;
		14'h3d18:	ff_dbi <= 8'h00;
		14'h3d19:	ff_dbi <= 8'h00;
		14'h3d1a:	ff_dbi <= 8'h00;
		14'h3d1b:	ff_dbi <= 8'h00;
		14'h3d1c:	ff_dbi <= 8'h00;
		14'h3d1d:	ff_dbi <= 8'h00;
		14'h3d1e:	ff_dbi <= 8'h00;
		14'h3d1f:	ff_dbi <= 8'h00;
		14'h3d20:	ff_dbi <= 8'h00;
		14'h3d21:	ff_dbi <= 8'h00;
		14'h3d22:	ff_dbi <= 8'h00;
		14'h3d23:	ff_dbi <= 8'h00;
		14'h3d24:	ff_dbi <= 8'h00;
		14'h3d25:	ff_dbi <= 8'h00;
		14'h3d26:	ff_dbi <= 8'h00;
		14'h3d27:	ff_dbi <= 8'h00;
		14'h3d28:	ff_dbi <= 8'h00;
		14'h3d29:	ff_dbi <= 8'h00;
		14'h3d2a:	ff_dbi <= 8'h00;
		14'h3d2b:	ff_dbi <= 8'h00;
		14'h3d2c:	ff_dbi <= 8'h00;
		14'h3d2d:	ff_dbi <= 8'h00;
		14'h3d2e:	ff_dbi <= 8'h00;
		14'h3d2f:	ff_dbi <= 8'h00;
		14'h3d30:	ff_dbi <= 8'h00;
		14'h3d31:	ff_dbi <= 8'h00;
		14'h3d32:	ff_dbi <= 8'h00;
		14'h3d33:	ff_dbi <= 8'h00;
		14'h3d34:	ff_dbi <= 8'h00;
		14'h3d35:	ff_dbi <= 8'h00;
		14'h3d36:	ff_dbi <= 8'h00;
		14'h3d37:	ff_dbi <= 8'h00;
		14'h3d38:	ff_dbi <= 8'h00;
		14'h3d39:	ff_dbi <= 8'h00;
		14'h3d3a:	ff_dbi <= 8'h00;
		14'h3d3b:	ff_dbi <= 8'h00;
		14'h3d3c:	ff_dbi <= 8'h00;
		14'h3d3d:	ff_dbi <= 8'h00;
		14'h3d3e:	ff_dbi <= 8'h00;
		14'h3d3f:	ff_dbi <= 8'h00;
		14'h3d40:	ff_dbi <= 8'h00;
		14'h3d41:	ff_dbi <= 8'h00;
		14'h3d42:	ff_dbi <= 8'h00;
		14'h3d43:	ff_dbi <= 8'h00;
		14'h3d44:	ff_dbi <= 8'h00;
		14'h3d45:	ff_dbi <= 8'h00;
		14'h3d46:	ff_dbi <= 8'h00;
		14'h3d47:	ff_dbi <= 8'h00;
		14'h3d48:	ff_dbi <= 8'h00;
		14'h3d49:	ff_dbi <= 8'h00;
		14'h3d4a:	ff_dbi <= 8'h00;
		14'h3d4b:	ff_dbi <= 8'h00;
		14'h3d4c:	ff_dbi <= 8'h00;
		14'h3d4d:	ff_dbi <= 8'h00;
		14'h3d4e:	ff_dbi <= 8'h00;
		14'h3d4f:	ff_dbi <= 8'h00;
		14'h3d50:	ff_dbi <= 8'h00;
		14'h3d51:	ff_dbi <= 8'h00;
		14'h3d52:	ff_dbi <= 8'h00;
		14'h3d53:	ff_dbi <= 8'h00;
		14'h3d54:	ff_dbi <= 8'h00;
		14'h3d55:	ff_dbi <= 8'h00;
		14'h3d56:	ff_dbi <= 8'h00;
		14'h3d57:	ff_dbi <= 8'h00;
		14'h3d58:	ff_dbi <= 8'h00;
		14'h3d59:	ff_dbi <= 8'h00;
		14'h3d5a:	ff_dbi <= 8'h00;
		14'h3d5b:	ff_dbi <= 8'h00;
		14'h3d5c:	ff_dbi <= 8'h00;
		14'h3d5d:	ff_dbi <= 8'h00;
		14'h3d5e:	ff_dbi <= 8'h00;
		14'h3d5f:	ff_dbi <= 8'h00;
		14'h3d60:	ff_dbi <= 8'h00;
		14'h3d61:	ff_dbi <= 8'h00;
		14'h3d62:	ff_dbi <= 8'h00;
		14'h3d63:	ff_dbi <= 8'h00;
		14'h3d64:	ff_dbi <= 8'h00;
		14'h3d65:	ff_dbi <= 8'h00;
		14'h3d66:	ff_dbi <= 8'h00;
		14'h3d67:	ff_dbi <= 8'h00;
		14'h3d68:	ff_dbi <= 8'h00;
		14'h3d69:	ff_dbi <= 8'h00;
		14'h3d6a:	ff_dbi <= 8'h00;
		14'h3d6b:	ff_dbi <= 8'h00;
		14'h3d6c:	ff_dbi <= 8'h00;
		14'h3d6d:	ff_dbi <= 8'h00;
		14'h3d6e:	ff_dbi <= 8'h00;
		14'h3d6f:	ff_dbi <= 8'h00;
		14'h3d70:	ff_dbi <= 8'h00;
		14'h3d71:	ff_dbi <= 8'h00;
		14'h3d72:	ff_dbi <= 8'h00;
		14'h3d73:	ff_dbi <= 8'h00;
		14'h3d74:	ff_dbi <= 8'h00;
		14'h3d75:	ff_dbi <= 8'h00;
		14'h3d76:	ff_dbi <= 8'h00;
		14'h3d77:	ff_dbi <= 8'h00;
		14'h3d78:	ff_dbi <= 8'h00;
		14'h3d79:	ff_dbi <= 8'h00;
		14'h3d7a:	ff_dbi <= 8'h00;
		14'h3d7b:	ff_dbi <= 8'h00;
		14'h3d7c:	ff_dbi <= 8'h00;
		14'h3d7d:	ff_dbi <= 8'h00;
		14'h3d7e:	ff_dbi <= 8'h00;
		14'h3d7f:	ff_dbi <= 8'h00;
		14'h3d80:	ff_dbi <= 8'h00;
		14'h3d81:	ff_dbi <= 8'h00;
		14'h3d82:	ff_dbi <= 8'h00;
		14'h3d83:	ff_dbi <= 8'h00;
		14'h3d84:	ff_dbi <= 8'h00;
		14'h3d85:	ff_dbi <= 8'h00;
		14'h3d86:	ff_dbi <= 8'h00;
		14'h3d87:	ff_dbi <= 8'h00;
		14'h3d88:	ff_dbi <= 8'h00;
		14'h3d89:	ff_dbi <= 8'h00;
		14'h3d8a:	ff_dbi <= 8'h00;
		14'h3d8b:	ff_dbi <= 8'h00;
		14'h3d8c:	ff_dbi <= 8'h00;
		14'h3d8d:	ff_dbi <= 8'h00;
		14'h3d8e:	ff_dbi <= 8'h00;
		14'h3d8f:	ff_dbi <= 8'h00;
		14'h3d90:	ff_dbi <= 8'h00;
		14'h3d91:	ff_dbi <= 8'h00;
		14'h3d92:	ff_dbi <= 8'h00;
		14'h3d93:	ff_dbi <= 8'h00;
		14'h3d94:	ff_dbi <= 8'h00;
		14'h3d95:	ff_dbi <= 8'h00;
		14'h3d96:	ff_dbi <= 8'h00;
		14'h3d97:	ff_dbi <= 8'h00;
		14'h3d98:	ff_dbi <= 8'h00;
		14'h3d99:	ff_dbi <= 8'h00;
		14'h3d9a:	ff_dbi <= 8'h00;
		14'h3d9b:	ff_dbi <= 8'h00;
		14'h3d9c:	ff_dbi <= 8'h00;
		14'h3d9d:	ff_dbi <= 8'h00;
		14'h3d9e:	ff_dbi <= 8'h00;
		14'h3d9f:	ff_dbi <= 8'h00;
		14'h3da0:	ff_dbi <= 8'h00;
		14'h3da1:	ff_dbi <= 8'h00;
		14'h3da2:	ff_dbi <= 8'h00;
		14'h3da3:	ff_dbi <= 8'h00;
		14'h3da4:	ff_dbi <= 8'h00;
		14'h3da5:	ff_dbi <= 8'h00;
		14'h3da6:	ff_dbi <= 8'h00;
		14'h3da7:	ff_dbi <= 8'h00;
		14'h3da8:	ff_dbi <= 8'h00;
		14'h3da9:	ff_dbi <= 8'h00;
		14'h3daa:	ff_dbi <= 8'h00;
		14'h3dab:	ff_dbi <= 8'h00;
		14'h3dac:	ff_dbi <= 8'h00;
		14'h3dad:	ff_dbi <= 8'h00;
		14'h3dae:	ff_dbi <= 8'h00;
		14'h3daf:	ff_dbi <= 8'h00;
		14'h3db0:	ff_dbi <= 8'h00;
		14'h3db1:	ff_dbi <= 8'h00;
		14'h3db2:	ff_dbi <= 8'h00;
		14'h3db3:	ff_dbi <= 8'h00;
		14'h3db4:	ff_dbi <= 8'h00;
		14'h3db5:	ff_dbi <= 8'h00;
		14'h3db6:	ff_dbi <= 8'h00;
		14'h3db7:	ff_dbi <= 8'h00;
		14'h3db8:	ff_dbi <= 8'h00;
		14'h3db9:	ff_dbi <= 8'h00;
		14'h3dba:	ff_dbi <= 8'h00;
		14'h3dbb:	ff_dbi <= 8'h00;
		14'h3dbc:	ff_dbi <= 8'h00;
		14'h3dbd:	ff_dbi <= 8'h00;
		14'h3dbe:	ff_dbi <= 8'h00;
		14'h3dbf:	ff_dbi <= 8'h00;
		14'h3dc0:	ff_dbi <= 8'h00;
		14'h3dc1:	ff_dbi <= 8'h00;
		14'h3dc2:	ff_dbi <= 8'h00;
		14'h3dc3:	ff_dbi <= 8'h00;
		14'h3dc4:	ff_dbi <= 8'h00;
		14'h3dc5:	ff_dbi <= 8'h00;
		14'h3dc6:	ff_dbi <= 8'h00;
		14'h3dc7:	ff_dbi <= 8'h00;
		14'h3dc8:	ff_dbi <= 8'h00;
		14'h3dc9:	ff_dbi <= 8'h00;
		14'h3dca:	ff_dbi <= 8'h00;
		14'h3dcb:	ff_dbi <= 8'h00;
		14'h3dcc:	ff_dbi <= 8'h00;
		14'h3dcd:	ff_dbi <= 8'h00;
		14'h3dce:	ff_dbi <= 8'h00;
		14'h3dcf:	ff_dbi <= 8'h00;
		14'h3dd0:	ff_dbi <= 8'h00;
		14'h3dd1:	ff_dbi <= 8'h00;
		14'h3dd2:	ff_dbi <= 8'h00;
		14'h3dd3:	ff_dbi <= 8'h00;
		14'h3dd4:	ff_dbi <= 8'h00;
		14'h3dd5:	ff_dbi <= 8'h00;
		14'h3dd6:	ff_dbi <= 8'h00;
		14'h3dd7:	ff_dbi <= 8'h00;
		14'h3dd8:	ff_dbi <= 8'h00;
		14'h3dd9:	ff_dbi <= 8'h00;
		14'h3dda:	ff_dbi <= 8'h00;
		14'h3ddb:	ff_dbi <= 8'h00;
		14'h3ddc:	ff_dbi <= 8'h00;
		14'h3ddd:	ff_dbi <= 8'h00;
		14'h3dde:	ff_dbi <= 8'h00;
		14'h3ddf:	ff_dbi <= 8'h00;
		14'h3de0:	ff_dbi <= 8'h00;
		14'h3de1:	ff_dbi <= 8'h00;
		14'h3de2:	ff_dbi <= 8'h00;
		14'h3de3:	ff_dbi <= 8'h00;
		14'h3de4:	ff_dbi <= 8'h00;
		14'h3de5:	ff_dbi <= 8'h00;
		14'h3de6:	ff_dbi <= 8'h00;
		14'h3de7:	ff_dbi <= 8'h00;
		14'h3de8:	ff_dbi <= 8'h00;
		14'h3de9:	ff_dbi <= 8'h00;
		14'h3dea:	ff_dbi <= 8'h00;
		14'h3deb:	ff_dbi <= 8'h00;
		14'h3dec:	ff_dbi <= 8'h00;
		14'h3ded:	ff_dbi <= 8'h00;
		14'h3dee:	ff_dbi <= 8'h00;
		14'h3def:	ff_dbi <= 8'h00;
		14'h3df0:	ff_dbi <= 8'h00;
		14'h3df1:	ff_dbi <= 8'h00;
		14'h3df2:	ff_dbi <= 8'h00;
		14'h3df3:	ff_dbi <= 8'h00;
		14'h3df4:	ff_dbi <= 8'h00;
		14'h3df5:	ff_dbi <= 8'h00;
		14'h3df6:	ff_dbi <= 8'h00;
		14'h3df7:	ff_dbi <= 8'h00;
		14'h3df8:	ff_dbi <= 8'h00;
		14'h3df9:	ff_dbi <= 8'h00;
		14'h3dfa:	ff_dbi <= 8'h00;
		14'h3dfb:	ff_dbi <= 8'h00;
		14'h3dfc:	ff_dbi <= 8'h00;
		14'h3dfd:	ff_dbi <= 8'h00;
		14'h3dfe:	ff_dbi <= 8'h00;
		14'h3dff:	ff_dbi <= 8'h00;
		14'h3e00:	ff_dbi <= 8'h00;
		14'h3e01:	ff_dbi <= 8'h00;
		14'h3e02:	ff_dbi <= 8'h00;
		14'h3e03:	ff_dbi <= 8'h00;
		14'h3e04:	ff_dbi <= 8'h00;
		14'h3e05:	ff_dbi <= 8'h00;
		14'h3e06:	ff_dbi <= 8'h00;
		14'h3e07:	ff_dbi <= 8'h00;
		14'h3e08:	ff_dbi <= 8'h00;
		14'h3e09:	ff_dbi <= 8'h00;
		14'h3e0a:	ff_dbi <= 8'h00;
		14'h3e0b:	ff_dbi <= 8'h00;
		14'h3e0c:	ff_dbi <= 8'h00;
		14'h3e0d:	ff_dbi <= 8'h00;
		14'h3e0e:	ff_dbi <= 8'h00;
		14'h3e0f:	ff_dbi <= 8'h00;
		14'h3e10:	ff_dbi <= 8'h00;
		14'h3e11:	ff_dbi <= 8'h00;
		14'h3e12:	ff_dbi <= 8'h00;
		14'h3e13:	ff_dbi <= 8'h00;
		14'h3e14:	ff_dbi <= 8'h00;
		14'h3e15:	ff_dbi <= 8'h00;
		14'h3e16:	ff_dbi <= 8'h00;
		14'h3e17:	ff_dbi <= 8'h00;
		14'h3e18:	ff_dbi <= 8'h00;
		14'h3e19:	ff_dbi <= 8'h00;
		14'h3e1a:	ff_dbi <= 8'h00;
		14'h3e1b:	ff_dbi <= 8'h00;
		14'h3e1c:	ff_dbi <= 8'h00;
		14'h3e1d:	ff_dbi <= 8'h00;
		14'h3e1e:	ff_dbi <= 8'h00;
		14'h3e1f:	ff_dbi <= 8'h00;
		14'h3e20:	ff_dbi <= 8'h00;
		14'h3e21:	ff_dbi <= 8'h00;
		14'h3e22:	ff_dbi <= 8'h00;
		14'h3e23:	ff_dbi <= 8'h00;
		14'h3e24:	ff_dbi <= 8'h00;
		14'h3e25:	ff_dbi <= 8'h00;
		14'h3e26:	ff_dbi <= 8'h00;
		14'h3e27:	ff_dbi <= 8'h00;
		14'h3e28:	ff_dbi <= 8'h00;
		14'h3e29:	ff_dbi <= 8'h00;
		14'h3e2a:	ff_dbi <= 8'h00;
		14'h3e2b:	ff_dbi <= 8'h00;
		14'h3e2c:	ff_dbi <= 8'h00;
		14'h3e2d:	ff_dbi <= 8'h00;
		14'h3e2e:	ff_dbi <= 8'h00;
		14'h3e2f:	ff_dbi <= 8'h00;
		14'h3e30:	ff_dbi <= 8'h00;
		14'h3e31:	ff_dbi <= 8'h00;
		14'h3e32:	ff_dbi <= 8'h00;
		14'h3e33:	ff_dbi <= 8'h00;
		14'h3e34:	ff_dbi <= 8'h00;
		14'h3e35:	ff_dbi <= 8'h00;
		14'h3e36:	ff_dbi <= 8'h00;
		14'h3e37:	ff_dbi <= 8'h00;
		14'h3e38:	ff_dbi <= 8'h00;
		14'h3e39:	ff_dbi <= 8'h00;
		14'h3e3a:	ff_dbi <= 8'h00;
		14'h3e3b:	ff_dbi <= 8'h00;
		14'h3e3c:	ff_dbi <= 8'h00;
		14'h3e3d:	ff_dbi <= 8'h00;
		14'h3e3e:	ff_dbi <= 8'h00;
		14'h3e3f:	ff_dbi <= 8'h00;
		14'h3e40:	ff_dbi <= 8'h00;
		14'h3e41:	ff_dbi <= 8'h00;
		14'h3e42:	ff_dbi <= 8'h00;
		14'h3e43:	ff_dbi <= 8'h00;
		14'h3e44:	ff_dbi <= 8'h00;
		14'h3e45:	ff_dbi <= 8'h00;
		14'h3e46:	ff_dbi <= 8'h00;
		14'h3e47:	ff_dbi <= 8'h00;
		14'h3e48:	ff_dbi <= 8'h00;
		14'h3e49:	ff_dbi <= 8'h00;
		14'h3e4a:	ff_dbi <= 8'h00;
		14'h3e4b:	ff_dbi <= 8'h00;
		14'h3e4c:	ff_dbi <= 8'h00;
		14'h3e4d:	ff_dbi <= 8'h00;
		14'h3e4e:	ff_dbi <= 8'h00;
		14'h3e4f:	ff_dbi <= 8'h00;
		14'h3e50:	ff_dbi <= 8'h00;
		14'h3e51:	ff_dbi <= 8'h00;
		14'h3e52:	ff_dbi <= 8'h00;
		14'h3e53:	ff_dbi <= 8'h00;
		14'h3e54:	ff_dbi <= 8'h00;
		14'h3e55:	ff_dbi <= 8'h00;
		14'h3e56:	ff_dbi <= 8'h00;
		14'h3e57:	ff_dbi <= 8'h00;
		14'h3e58:	ff_dbi <= 8'h00;
		14'h3e59:	ff_dbi <= 8'h00;
		14'h3e5a:	ff_dbi <= 8'h00;
		14'h3e5b:	ff_dbi <= 8'h00;
		14'h3e5c:	ff_dbi <= 8'h00;
		14'h3e5d:	ff_dbi <= 8'h00;
		14'h3e5e:	ff_dbi <= 8'h00;
		14'h3e5f:	ff_dbi <= 8'h00;
		14'h3e60:	ff_dbi <= 8'h00;
		14'h3e61:	ff_dbi <= 8'h00;
		14'h3e62:	ff_dbi <= 8'h00;
		14'h3e63:	ff_dbi <= 8'h00;
		14'h3e64:	ff_dbi <= 8'h00;
		14'h3e65:	ff_dbi <= 8'h00;
		14'h3e66:	ff_dbi <= 8'h00;
		14'h3e67:	ff_dbi <= 8'h00;
		14'h3e68:	ff_dbi <= 8'h00;
		14'h3e69:	ff_dbi <= 8'h00;
		14'h3e6a:	ff_dbi <= 8'h00;
		14'h3e6b:	ff_dbi <= 8'h00;
		14'h3e6c:	ff_dbi <= 8'h00;
		14'h3e6d:	ff_dbi <= 8'h00;
		14'h3e6e:	ff_dbi <= 8'h00;
		14'h3e6f:	ff_dbi <= 8'h00;
		14'h3e70:	ff_dbi <= 8'h00;
		14'h3e71:	ff_dbi <= 8'h00;
		14'h3e72:	ff_dbi <= 8'h00;
		14'h3e73:	ff_dbi <= 8'h00;
		14'h3e74:	ff_dbi <= 8'h00;
		14'h3e75:	ff_dbi <= 8'h00;
		14'h3e76:	ff_dbi <= 8'h00;
		14'h3e77:	ff_dbi <= 8'h00;
		14'h3e78:	ff_dbi <= 8'h00;
		14'h3e79:	ff_dbi <= 8'h00;
		14'h3e7a:	ff_dbi <= 8'h00;
		14'h3e7b:	ff_dbi <= 8'h00;
		14'h3e7c:	ff_dbi <= 8'h00;
		14'h3e7d:	ff_dbi <= 8'h00;
		14'h3e7e:	ff_dbi <= 8'h00;
		14'h3e7f:	ff_dbi <= 8'h00;
		14'h3e80:	ff_dbi <= 8'h00;
		14'h3e81:	ff_dbi <= 8'h00;
		14'h3e82:	ff_dbi <= 8'h00;
		14'h3e83:	ff_dbi <= 8'h00;
		14'h3e84:	ff_dbi <= 8'h00;
		14'h3e85:	ff_dbi <= 8'h00;
		14'h3e86:	ff_dbi <= 8'h00;
		14'h3e87:	ff_dbi <= 8'h00;
		14'h3e88:	ff_dbi <= 8'h00;
		14'h3e89:	ff_dbi <= 8'h00;
		14'h3e8a:	ff_dbi <= 8'h00;
		14'h3e8b:	ff_dbi <= 8'h00;
		14'h3e8c:	ff_dbi <= 8'h00;
		14'h3e8d:	ff_dbi <= 8'h00;
		14'h3e8e:	ff_dbi <= 8'h00;
		14'h3e8f:	ff_dbi <= 8'h00;
		14'h3e90:	ff_dbi <= 8'h00;
		14'h3e91:	ff_dbi <= 8'h00;
		14'h3e92:	ff_dbi <= 8'h00;
		14'h3e93:	ff_dbi <= 8'h00;
		14'h3e94:	ff_dbi <= 8'h00;
		14'h3e95:	ff_dbi <= 8'h00;
		14'h3e96:	ff_dbi <= 8'h00;
		14'h3e97:	ff_dbi <= 8'h00;
		14'h3e98:	ff_dbi <= 8'h00;
		14'h3e99:	ff_dbi <= 8'h00;
		14'h3e9a:	ff_dbi <= 8'h00;
		14'h3e9b:	ff_dbi <= 8'h00;
		14'h3e9c:	ff_dbi <= 8'h00;
		14'h3e9d:	ff_dbi <= 8'h00;
		14'h3e9e:	ff_dbi <= 8'h00;
		14'h3e9f:	ff_dbi <= 8'h00;
		14'h3ea0:	ff_dbi <= 8'h00;
		14'h3ea1:	ff_dbi <= 8'h00;
		14'h3ea2:	ff_dbi <= 8'h00;
		14'h3ea3:	ff_dbi <= 8'h00;
		14'h3ea4:	ff_dbi <= 8'h00;
		14'h3ea5:	ff_dbi <= 8'h00;
		14'h3ea6:	ff_dbi <= 8'h00;
		14'h3ea7:	ff_dbi <= 8'h00;
		14'h3ea8:	ff_dbi <= 8'h00;
		14'h3ea9:	ff_dbi <= 8'h00;
		14'h3eaa:	ff_dbi <= 8'h00;
		14'h3eab:	ff_dbi <= 8'h00;
		14'h3eac:	ff_dbi <= 8'h00;
		14'h3ead:	ff_dbi <= 8'h00;
		14'h3eae:	ff_dbi <= 8'h00;
		14'h3eaf:	ff_dbi <= 8'h00;
		14'h3eb0:	ff_dbi <= 8'h00;
		14'h3eb1:	ff_dbi <= 8'h00;
		14'h3eb2:	ff_dbi <= 8'h00;
		14'h3eb3:	ff_dbi <= 8'h00;
		14'h3eb4:	ff_dbi <= 8'h00;
		14'h3eb5:	ff_dbi <= 8'h00;
		14'h3eb6:	ff_dbi <= 8'h00;
		14'h3eb7:	ff_dbi <= 8'h00;
		14'h3eb8:	ff_dbi <= 8'h00;
		14'h3eb9:	ff_dbi <= 8'h00;
		14'h3eba:	ff_dbi <= 8'h00;
		14'h3ebb:	ff_dbi <= 8'h00;
		14'h3ebc:	ff_dbi <= 8'h00;
		14'h3ebd:	ff_dbi <= 8'h00;
		14'h3ebe:	ff_dbi <= 8'h00;
		14'h3ebf:	ff_dbi <= 8'h00;
		14'h3ec0:	ff_dbi <= 8'h00;
		14'h3ec1:	ff_dbi <= 8'h00;
		14'h3ec2:	ff_dbi <= 8'h00;
		14'h3ec3:	ff_dbi <= 8'h00;
		14'h3ec4:	ff_dbi <= 8'h00;
		14'h3ec5:	ff_dbi <= 8'h00;
		14'h3ec6:	ff_dbi <= 8'h00;
		14'h3ec7:	ff_dbi <= 8'h00;
		14'h3ec8:	ff_dbi <= 8'h00;
		14'h3ec9:	ff_dbi <= 8'h00;
		14'h3eca:	ff_dbi <= 8'h00;
		14'h3ecb:	ff_dbi <= 8'h00;
		14'h3ecc:	ff_dbi <= 8'h00;
		14'h3ecd:	ff_dbi <= 8'h00;
		14'h3ece:	ff_dbi <= 8'h00;
		14'h3ecf:	ff_dbi <= 8'h00;
		14'h3ed0:	ff_dbi <= 8'h00;
		14'h3ed1:	ff_dbi <= 8'h00;
		14'h3ed2:	ff_dbi <= 8'h00;
		14'h3ed3:	ff_dbi <= 8'h00;
		14'h3ed4:	ff_dbi <= 8'h00;
		14'h3ed5:	ff_dbi <= 8'h00;
		14'h3ed6:	ff_dbi <= 8'h00;
		14'h3ed7:	ff_dbi <= 8'h00;
		14'h3ed8:	ff_dbi <= 8'h00;
		14'h3ed9:	ff_dbi <= 8'h00;
		14'h3eda:	ff_dbi <= 8'h00;
		14'h3edb:	ff_dbi <= 8'h00;
		14'h3edc:	ff_dbi <= 8'h00;
		14'h3edd:	ff_dbi <= 8'h00;
		14'h3ede:	ff_dbi <= 8'h00;
		14'h3edf:	ff_dbi <= 8'h00;
		14'h3ee0:	ff_dbi <= 8'h00;
		14'h3ee1:	ff_dbi <= 8'h00;
		14'h3ee2:	ff_dbi <= 8'h00;
		14'h3ee3:	ff_dbi <= 8'h00;
		14'h3ee4:	ff_dbi <= 8'h00;
		14'h3ee5:	ff_dbi <= 8'h00;
		14'h3ee6:	ff_dbi <= 8'h00;
		14'h3ee7:	ff_dbi <= 8'h00;
		14'h3ee8:	ff_dbi <= 8'h00;
		14'h3ee9:	ff_dbi <= 8'h00;
		14'h3eea:	ff_dbi <= 8'h00;
		14'h3eeb:	ff_dbi <= 8'h00;
		14'h3eec:	ff_dbi <= 8'h00;
		14'h3eed:	ff_dbi <= 8'h00;
		14'h3eee:	ff_dbi <= 8'h00;
		14'h3eef:	ff_dbi <= 8'h00;
		14'h3ef0:	ff_dbi <= 8'h00;
		14'h3ef1:	ff_dbi <= 8'h00;
		14'h3ef2:	ff_dbi <= 8'h00;
		14'h3ef3:	ff_dbi <= 8'h00;
		14'h3ef4:	ff_dbi <= 8'h00;
		14'h3ef5:	ff_dbi <= 8'h00;
		14'h3ef6:	ff_dbi <= 8'h00;
		14'h3ef7:	ff_dbi <= 8'h00;
		14'h3ef8:	ff_dbi <= 8'h00;
		14'h3ef9:	ff_dbi <= 8'h00;
		14'h3efa:	ff_dbi <= 8'h00;
		14'h3efb:	ff_dbi <= 8'h00;
		14'h3efc:	ff_dbi <= 8'h00;
		14'h3efd:	ff_dbi <= 8'h00;
		14'h3efe:	ff_dbi <= 8'h00;
		14'h3eff:	ff_dbi <= 8'h00;
		14'h3f00:	ff_dbi <= 8'h00;
		14'h3f01:	ff_dbi <= 8'h00;
		14'h3f02:	ff_dbi <= 8'h00;
		14'h3f03:	ff_dbi <= 8'h00;
		14'h3f04:	ff_dbi <= 8'h00;
		14'h3f05:	ff_dbi <= 8'h00;
		14'h3f06:	ff_dbi <= 8'h00;
		14'h3f07:	ff_dbi <= 8'h00;
		14'h3f08:	ff_dbi <= 8'h00;
		14'h3f09:	ff_dbi <= 8'h00;
		14'h3f0a:	ff_dbi <= 8'h00;
		14'h3f0b:	ff_dbi <= 8'h00;
		14'h3f0c:	ff_dbi <= 8'h00;
		14'h3f0d:	ff_dbi <= 8'h00;
		14'h3f0e:	ff_dbi <= 8'h00;
		14'h3f0f:	ff_dbi <= 8'h00;
		14'h3f10:	ff_dbi <= 8'h00;
		14'h3f11:	ff_dbi <= 8'h00;
		14'h3f12:	ff_dbi <= 8'h00;
		14'h3f13:	ff_dbi <= 8'h00;
		14'h3f14:	ff_dbi <= 8'h00;
		14'h3f15:	ff_dbi <= 8'h00;
		14'h3f16:	ff_dbi <= 8'h00;
		14'h3f17:	ff_dbi <= 8'h00;
		14'h3f18:	ff_dbi <= 8'h00;
		14'h3f19:	ff_dbi <= 8'h00;
		14'h3f1a:	ff_dbi <= 8'h00;
		14'h3f1b:	ff_dbi <= 8'h00;
		14'h3f1c:	ff_dbi <= 8'h00;
		14'h3f1d:	ff_dbi <= 8'h00;
		14'h3f1e:	ff_dbi <= 8'h00;
		14'h3f1f:	ff_dbi <= 8'h00;
		14'h3f20:	ff_dbi <= 8'h00;
		14'h3f21:	ff_dbi <= 8'h00;
		14'h3f22:	ff_dbi <= 8'h00;
		14'h3f23:	ff_dbi <= 8'h00;
		14'h3f24:	ff_dbi <= 8'h00;
		14'h3f25:	ff_dbi <= 8'h00;
		14'h3f26:	ff_dbi <= 8'h00;
		14'h3f27:	ff_dbi <= 8'h00;
		14'h3f28:	ff_dbi <= 8'h00;
		14'h3f29:	ff_dbi <= 8'h00;
		14'h3f2a:	ff_dbi <= 8'h00;
		14'h3f2b:	ff_dbi <= 8'h00;
		14'h3f2c:	ff_dbi <= 8'h00;
		14'h3f2d:	ff_dbi <= 8'h00;
		14'h3f2e:	ff_dbi <= 8'h00;
		14'h3f2f:	ff_dbi <= 8'h00;
		14'h3f30:	ff_dbi <= 8'h00;
		14'h3f31:	ff_dbi <= 8'h00;
		14'h3f32:	ff_dbi <= 8'h00;
		14'h3f33:	ff_dbi <= 8'h00;
		14'h3f34:	ff_dbi <= 8'h00;
		14'h3f35:	ff_dbi <= 8'h00;
		14'h3f36:	ff_dbi <= 8'h00;
		14'h3f37:	ff_dbi <= 8'h00;
		14'h3f38:	ff_dbi <= 8'h00;
		14'h3f39:	ff_dbi <= 8'h00;
		14'h3f3a:	ff_dbi <= 8'h00;
		14'h3f3b:	ff_dbi <= 8'h00;
		14'h3f3c:	ff_dbi <= 8'h00;
		14'h3f3d:	ff_dbi <= 8'h00;
		14'h3f3e:	ff_dbi <= 8'h00;
		14'h3f3f:	ff_dbi <= 8'h00;
		14'h3f40:	ff_dbi <= 8'h00;
		14'h3f41:	ff_dbi <= 8'h00;
		14'h3f42:	ff_dbi <= 8'h00;
		14'h3f43:	ff_dbi <= 8'h00;
		14'h3f44:	ff_dbi <= 8'h00;
		14'h3f45:	ff_dbi <= 8'h00;
		14'h3f46:	ff_dbi <= 8'h00;
		14'h3f47:	ff_dbi <= 8'h00;
		14'h3f48:	ff_dbi <= 8'h00;
		14'h3f49:	ff_dbi <= 8'h00;
		14'h3f4a:	ff_dbi <= 8'h00;
		14'h3f4b:	ff_dbi <= 8'h00;
		14'h3f4c:	ff_dbi <= 8'h00;
		14'h3f4d:	ff_dbi <= 8'h00;
		14'h3f4e:	ff_dbi <= 8'h00;
		14'h3f4f:	ff_dbi <= 8'h00;
		14'h3f50:	ff_dbi <= 8'h00;
		14'h3f51:	ff_dbi <= 8'h00;
		14'h3f52:	ff_dbi <= 8'h00;
		14'h3f53:	ff_dbi <= 8'h00;
		14'h3f54:	ff_dbi <= 8'h00;
		14'h3f55:	ff_dbi <= 8'h00;
		14'h3f56:	ff_dbi <= 8'h00;
		14'h3f57:	ff_dbi <= 8'h00;
		14'h3f58:	ff_dbi <= 8'h00;
		14'h3f59:	ff_dbi <= 8'h00;
		14'h3f5a:	ff_dbi <= 8'h00;
		14'h3f5b:	ff_dbi <= 8'h00;
		14'h3f5c:	ff_dbi <= 8'h00;
		14'h3f5d:	ff_dbi <= 8'h00;
		14'h3f5e:	ff_dbi <= 8'h00;
		14'h3f5f:	ff_dbi <= 8'h00;
		14'h3f60:	ff_dbi <= 8'h00;
		14'h3f61:	ff_dbi <= 8'h00;
		14'h3f62:	ff_dbi <= 8'h00;
		14'h3f63:	ff_dbi <= 8'h00;
		14'h3f64:	ff_dbi <= 8'h00;
		14'h3f65:	ff_dbi <= 8'h00;
		14'h3f66:	ff_dbi <= 8'h00;
		14'h3f67:	ff_dbi <= 8'h00;
		14'h3f68:	ff_dbi <= 8'h00;
		14'h3f69:	ff_dbi <= 8'h00;
		14'h3f6a:	ff_dbi <= 8'h00;
		14'h3f6b:	ff_dbi <= 8'h00;
		14'h3f6c:	ff_dbi <= 8'h00;
		14'h3f6d:	ff_dbi <= 8'h00;
		14'h3f6e:	ff_dbi <= 8'h00;
		14'h3f6f:	ff_dbi <= 8'h00;
		14'h3f70:	ff_dbi <= 8'h00;
		14'h3f71:	ff_dbi <= 8'h00;
		14'h3f72:	ff_dbi <= 8'h00;
		14'h3f73:	ff_dbi <= 8'h00;
		14'h3f74:	ff_dbi <= 8'h00;
		14'h3f75:	ff_dbi <= 8'h00;
		14'h3f76:	ff_dbi <= 8'h00;
		14'h3f77:	ff_dbi <= 8'h00;
		14'h3f78:	ff_dbi <= 8'h00;
		14'h3f79:	ff_dbi <= 8'h00;
		14'h3f7a:	ff_dbi <= 8'h00;
		14'h3f7b:	ff_dbi <= 8'h00;
		14'h3f7c:	ff_dbi <= 8'h00;
		14'h3f7d:	ff_dbi <= 8'h00;
		14'h3f7e:	ff_dbi <= 8'h00;
		14'h3f7f:	ff_dbi <= 8'h00;
		14'h3f80:	ff_dbi <= 8'h00;
		14'h3f81:	ff_dbi <= 8'h00;
		14'h3f82:	ff_dbi <= 8'h00;
		14'h3f83:	ff_dbi <= 8'h00;
		14'h3f84:	ff_dbi <= 8'h00;
		14'h3f85:	ff_dbi <= 8'h00;
		14'h3f86:	ff_dbi <= 8'h00;
		14'h3f87:	ff_dbi <= 8'h00;
		14'h3f88:	ff_dbi <= 8'h00;
		14'h3f89:	ff_dbi <= 8'h00;
		14'h3f8a:	ff_dbi <= 8'h00;
		14'h3f8b:	ff_dbi <= 8'h00;
		14'h3f8c:	ff_dbi <= 8'h00;
		14'h3f8d:	ff_dbi <= 8'h00;
		14'h3f8e:	ff_dbi <= 8'h00;
		14'h3f8f:	ff_dbi <= 8'h00;
		14'h3f90:	ff_dbi <= 8'h00;
		14'h3f91:	ff_dbi <= 8'h00;
		14'h3f92:	ff_dbi <= 8'h00;
		14'h3f93:	ff_dbi <= 8'h00;
		14'h3f94:	ff_dbi <= 8'h00;
		14'h3f95:	ff_dbi <= 8'h00;
		14'h3f96:	ff_dbi <= 8'h00;
		14'h3f97:	ff_dbi <= 8'h00;
		14'h3f98:	ff_dbi <= 8'h00;
		14'h3f99:	ff_dbi <= 8'h00;
		14'h3f9a:	ff_dbi <= 8'h00;
		14'h3f9b:	ff_dbi <= 8'h00;
		14'h3f9c:	ff_dbi <= 8'h00;
		14'h3f9d:	ff_dbi <= 8'h00;
		14'h3f9e:	ff_dbi <= 8'h00;
		14'h3f9f:	ff_dbi <= 8'h00;
		14'h3fa0:	ff_dbi <= 8'h00;
		14'h3fa1:	ff_dbi <= 8'h00;
		14'h3fa2:	ff_dbi <= 8'h00;
		14'h3fa3:	ff_dbi <= 8'h00;
		14'h3fa4:	ff_dbi <= 8'h00;
		14'h3fa5:	ff_dbi <= 8'h00;
		14'h3fa6:	ff_dbi <= 8'h00;
		14'h3fa7:	ff_dbi <= 8'h00;
		14'h3fa8:	ff_dbi <= 8'h00;
		14'h3fa9:	ff_dbi <= 8'h00;
		14'h3faa:	ff_dbi <= 8'h00;
		14'h3fab:	ff_dbi <= 8'h00;
		14'h3fac:	ff_dbi <= 8'h00;
		14'h3fad:	ff_dbi <= 8'h00;
		14'h3fae:	ff_dbi <= 8'h00;
		14'h3faf:	ff_dbi <= 8'h00;
		14'h3fb0:	ff_dbi <= 8'h00;
		14'h3fb1:	ff_dbi <= 8'h00;
		14'h3fb2:	ff_dbi <= 8'h00;
		14'h3fb3:	ff_dbi <= 8'h00;
		14'h3fb4:	ff_dbi <= 8'h00;
		14'h3fb5:	ff_dbi <= 8'h00;
		14'h3fb6:	ff_dbi <= 8'h00;
		14'h3fb7:	ff_dbi <= 8'h00;
		14'h3fb8:	ff_dbi <= 8'h00;
		14'h3fb9:	ff_dbi <= 8'h00;
		14'h3fba:	ff_dbi <= 8'h00;
		14'h3fbb:	ff_dbi <= 8'h00;
		14'h3fbc:	ff_dbi <= 8'h00;
		14'h3fbd:	ff_dbi <= 8'h00;
		14'h3fbe:	ff_dbi <= 8'h00;
		14'h3fbf:	ff_dbi <= 8'h00;
		14'h3fc0:	ff_dbi <= 8'h00;
		14'h3fc1:	ff_dbi <= 8'h00;
		14'h3fc2:	ff_dbi <= 8'h00;
		14'h3fc3:	ff_dbi <= 8'h00;
		14'h3fc4:	ff_dbi <= 8'h00;
		14'h3fc5:	ff_dbi <= 8'h00;
		14'h3fc6:	ff_dbi <= 8'h00;
		14'h3fc7:	ff_dbi <= 8'h00;
		14'h3fc8:	ff_dbi <= 8'h00;
		14'h3fc9:	ff_dbi <= 8'h00;
		14'h3fca:	ff_dbi <= 8'h00;
		14'h3fcb:	ff_dbi <= 8'h00;
		14'h3fcc:	ff_dbi <= 8'h00;
		14'h3fcd:	ff_dbi <= 8'h00;
		14'h3fce:	ff_dbi <= 8'h00;
		14'h3fcf:	ff_dbi <= 8'h00;
		14'h3fd0:	ff_dbi <= 8'h00;
		14'h3fd1:	ff_dbi <= 8'h00;
		14'h3fd2:	ff_dbi <= 8'h00;
		14'h3fd3:	ff_dbi <= 8'h00;
		14'h3fd4:	ff_dbi <= 8'h00;
		14'h3fd5:	ff_dbi <= 8'h00;
		14'h3fd6:	ff_dbi <= 8'h00;
		14'h3fd7:	ff_dbi <= 8'h00;
		14'h3fd8:	ff_dbi <= 8'h00;
		14'h3fd9:	ff_dbi <= 8'h00;
		14'h3fda:	ff_dbi <= 8'h00;
		14'h3fdb:	ff_dbi <= 8'h00;
		14'h3fdc:	ff_dbi <= 8'h00;
		14'h3fdd:	ff_dbi <= 8'h00;
		14'h3fde:	ff_dbi <= 8'h00;
		14'h3fdf:	ff_dbi <= 8'h00;
		14'h3fe0:	ff_dbi <= 8'h00;
		14'h3fe1:	ff_dbi <= 8'h00;
		14'h3fe2:	ff_dbi <= 8'h00;
		14'h3fe3:	ff_dbi <= 8'h00;
		14'h3fe4:	ff_dbi <= 8'h00;
		14'h3fe5:	ff_dbi <= 8'h00;
		14'h3fe6:	ff_dbi <= 8'h00;
		14'h3fe7:	ff_dbi <= 8'h00;
		14'h3fe8:	ff_dbi <= 8'h00;
		14'h3fe9:	ff_dbi <= 8'h00;
		14'h3fea:	ff_dbi <= 8'h00;
		14'h3feb:	ff_dbi <= 8'h00;
		14'h3fec:	ff_dbi <= 8'h00;
		14'h3fed:	ff_dbi <= 8'h00;
		14'h3fee:	ff_dbi <= 8'h00;
		14'h3fef:	ff_dbi <= 8'h00;
		14'h3ff0:	ff_dbi <= 8'h00;
		14'h3ff1:	ff_dbi <= 8'h00;
		14'h3ff2:	ff_dbi <= 8'h00;
		14'h3ff3:	ff_dbi <= 8'h00;
		14'h3ff4:	ff_dbi <= 8'h00;
		14'h3ff5:	ff_dbi <= 8'h00;
		14'h3ff6:	ff_dbi <= 8'h00;
		14'h3ff7:	ff_dbi <= 8'h00;
		14'h3ff8:	ff_dbi <= 8'h00;
		14'h3ff9:	ff_dbi <= 8'h00;
		14'h3ffa:	ff_dbi <= 8'h00;
		14'h3ffb:	ff_dbi <= 8'h00;
		14'h3ffc:	ff_dbi <= 8'h00;
		14'h3ffd:	ff_dbi <= 8'h00;
		14'h3ffe:	ff_dbi <= 8'h00;
		14'h3fff:	ff_dbi <= 8'h00;
		default:	ff_dbi <= 8'hxx;
		endcase
	end
endmodule
