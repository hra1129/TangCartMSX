parameter PLL_FCLKIN = "50";
parameter CLK_PERIOD = 20;
parameter SSC_DIR = 1'b0;
parameter SSC_EN = "TRUE";
parameter FRAC_DIV = 31'h1008AEFB; 
parameter PLL_ODIV0 = 8'd112;
parameter PLL_IDIV = 7'd1;
parameter PLL_FBDIV = 7'd1;
parameter SSC_CLKDIV = 28'd1516;
parameter SSC_STEP = 31'd3551;
