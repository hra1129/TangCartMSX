// --------------------------------------------------------------------
// IP_MSXMUSIC_ROM
// --------------------------------------------------------------------

module ip_msxmusic_rom (
	input			clk,
	input			n_cs,
	input			n_rd,
	input	[13:0]	address,
	output	[7:0]	rdata,
	output			rdata_en
);
	reg		[7:0]	ff_rdata;
	reg				ff_rdata_en;

	always @( posedge clk ) begin
		if( !n_cs && !n_rd ) begin
			case( address )
			14'd0: ff_rdata <= 8'h41;
			14'd1: ff_rdata <= 8'h42;
			14'd2: ff_rdata <= 8'h00;
			14'd3: ff_rdata <= 8'h00;
			14'd4: ff_rdata <= 8'h82;
			14'd5: ff_rdata <= 8'h40;
			14'd6: ff_rdata <= 8'h00;
			14'd7: ff_rdata <= 8'h00;
			14'd8: ff_rdata <= 8'h00;
			14'd9: ff_rdata <= 8'h00;
			14'd10: ff_rdata <= 8'h00;
			14'd11: ff_rdata <= 8'h00;
			14'd12: ff_rdata <= 8'h00;
			14'd13: ff_rdata <= 8'h00;
			14'd14: ff_rdata <= 8'h00;
			14'd15: ff_rdata <= 8'h00;
			14'd16: ff_rdata <= 8'h00;
			14'd17: ff_rdata <= 8'h00;
			14'd18: ff_rdata <= 8'h00;
			14'd19: ff_rdata <= 8'h00;
			14'd20: ff_rdata <= 8'h00;
			14'd21: ff_rdata <= 8'h00;
			14'd22: ff_rdata <= 8'h00;
			14'd23: ff_rdata <= 8'h00;
			14'd24: ff_rdata <= 8'h50;
			14'd25: ff_rdata <= 8'h41;
			14'd26: ff_rdata <= 8'h43;
			14'd27: ff_rdata <= 8'h32;
			14'd28: ff_rdata <= 8'h4F;
			14'd29: ff_rdata <= 8'h50;
			14'd30: ff_rdata <= 8'h4C;
			14'd31: ff_rdata <= 8'h4C;
			14'd32: ff_rdata <= 8'hC3;
			14'd33: ff_rdata <= 8'h64;
			14'd34: ff_rdata <= 8'h40;
			14'd35: ff_rdata <= 8'hC3;
			14'd36: ff_rdata <= 8'h5E;
			14'd37: ff_rdata <= 8'h40;
			14'd38: ff_rdata <= 8'hC3;
			14'd39: ff_rdata <= 8'h48;
			14'd40: ff_rdata <= 8'h40;
			14'd41: ff_rdata <= 8'hC3;
			14'd42: ff_rdata <= 8'h2F;
			14'd43: ff_rdata <= 8'h40;
			14'd44: ff_rdata <= 8'hC3;
			14'd45: ff_rdata <= 8'h3D;
			14'd46: ff_rdata <= 8'h40;
			14'd47: ff_rdata <= 8'hC5;
			14'd48: ff_rdata <= 8'h01;
			14'd49: ff_rdata <= 8'hF7;
			14'd50: ff_rdata <= 8'h7F;
			14'd51: ff_rdata <= 8'h0A;
			14'd52: ff_rdata <= 8'h08;
			14'd53: ff_rdata <= 8'h7B;
			14'd54: ff_rdata <= 8'h02;
			14'd55: ff_rdata <= 8'h7E;
			14'd56: ff_rdata <= 8'h08;
			14'd57: ff_rdata <= 8'h02;
			14'd58: ff_rdata <= 8'h08;
			14'd59: ff_rdata <= 8'hC1;
			14'd60: ff_rdata <= 8'hC9;
			14'd61: ff_rdata <= 8'hCD;
			14'd62: ff_rdata <= 8'h2F;
			14'd63: ff_rdata <= 8'h40;
			14'd64: ff_rdata <= 8'h57;
			14'd65: ff_rdata <= 8'h23;
			14'd66: ff_rdata <= 8'hCD;
			14'd67: ff_rdata <= 8'h2F;
			14'd68: ff_rdata <= 8'h40;
			14'd69: ff_rdata <= 8'h67;
			14'd70: ff_rdata <= 8'h6A;
			14'd71: ff_rdata <= 8'hC9;
			14'd72: ff_rdata <= 8'h3A;
			14'd73: ff_rdata <= 8'hF7;
			14'd74: ff_rdata <= 8'h7F;
			14'd75: ff_rdata <= 8'h08;
			14'd76: ff_rdata <= 8'hD9;
			14'd77: ff_rdata <= 8'hE1;
			14'd78: ff_rdata <= 8'hD1;
			14'd79: ff_rdata <= 8'hD5;
			14'd80: ff_rdata <= 8'hE5;
			14'd81: ff_rdata <= 8'h7B;
			14'd82: ff_rdata <= 8'hD9;
			14'd83: ff_rdata <= 8'h32;
			14'd84: ff_rdata <= 8'hF7;
			14'd85: ff_rdata <= 8'h7F;
			14'd86: ff_rdata <= 8'hEB;
			14'd87: ff_rdata <= 8'hED;
			14'd88: ff_rdata <= 8'hB0;
			14'd89: ff_rdata <= 8'h08;
			14'd90: ff_rdata <= 8'h32;
			14'd91: ff_rdata <= 8'hF7;
			14'd92: ff_rdata <= 8'h7F;
			14'd93: ff_rdata <= 8'hC9;
			14'd94: ff_rdata <= 8'hC5;
			14'd95: ff_rdata <= 8'hD9;
			14'd96: ff_rdata <= 8'hE1;
			14'd97: ff_rdata <= 8'hC3;
			14'd98: ff_rdata <= 8'h64;
			14'd99: ff_rdata <= 8'h40;
			14'd100: ff_rdata <= 8'hD9;
			14'd101: ff_rdata <= 8'h08;
			14'd102: ff_rdata <= 8'h3A;
			14'd103: ff_rdata <= 8'hF7;
			14'd104: ff_rdata <= 8'h7F;
			14'd105: ff_rdata <= 8'hF5;
			14'd106: ff_rdata <= 8'h7B;
			14'd107: ff_rdata <= 8'h32;
			14'd108: ff_rdata <= 8'hF7;
			14'd109: ff_rdata <= 8'h7F;
			14'd110: ff_rdata <= 8'h11;
			14'd111: ff_rdata <= 8'h76;
			14'd112: ff_rdata <= 8'h40;
			14'd113: ff_rdata <= 8'hD5;
			14'd114: ff_rdata <= 8'hE5;
			14'd115: ff_rdata <= 8'h08;
			14'd116: ff_rdata <= 8'hD9;
			14'd117: ff_rdata <= 8'hC9;
			14'd118: ff_rdata <= 8'h08;
			14'd119: ff_rdata <= 8'hF1;
			14'd120: ff_rdata <= 8'h32;
			14'd121: ff_rdata <= 8'hF7;
			14'd122: ff_rdata <= 8'h7F;
			14'd123: ff_rdata <= 8'h08;
			14'd124: ff_rdata <= 8'hC9;
			14'd125: ff_rdata <= 8'h00;
			14'd126: ff_rdata <= 8'h00;
			14'd127: ff_rdata <= 8'h00;
			14'd128: ff_rdata <= 8'h00;
			14'd129: ff_rdata <= 8'h50;
			14'd130: ff_rdata <= 8'hE5;
			14'd131: ff_rdata <= 8'h21;
			14'd132: ff_rdata <= 8'h89;
			14'd133: ff_rdata <= 8'hFD;
			14'd134: ff_rdata <= 8'h11;
			14'd135: ff_rdata <= 8'hB3;
			14'd136: ff_rdata <= 8'h40;
			14'd137: ff_rdata <= 8'h1A;
			14'd138: ff_rdata <= 8'hBE;
			14'd139: ff_rdata <= 8'h23;
			14'd140: ff_rdata <= 8'h13;
			14'd141: ff_rdata <= 8'h20;
			14'd142: ff_rdata <= 8'h17;
			14'd143: ff_rdata <= 8'hA7;
			14'd144: ff_rdata <= 8'h20;
			14'd145: ff_rdata <= 8'hF7;
			14'd146: ff_rdata <= 8'hE1;
			14'd147: ff_rdata <= 8'h3A;
			14'd148: ff_rdata <= 8'h06;
			14'd149: ff_rdata <= 8'h50;
			14'd150: ff_rdata <= 8'h3C;
			14'd151: ff_rdata <= 8'hC4;
			14'd152: ff_rdata <= 8'h06;
			14'd153: ff_rdata <= 8'h50;
			14'd154: ff_rdata <= 8'h1E;
			14'd155: ff_rdata <= 8'h01;
			14'd156: ff_rdata <= 8'h21;
			14'd157: ff_rdata <= 8'h80;
			14'd158: ff_rdata <= 8'h40;
			14'd159: ff_rdata <= 8'hCD;
			14'd160: ff_rdata <= 8'h2C;
			14'd161: ff_rdata <= 8'h40;
			14'd162: ff_rdata <= 8'hD9;
			14'd163: ff_rdata <= 8'hC3;
			14'd164: ff_rdata <= 8'h20;
			14'd165: ff_rdata <= 8'h40;
			14'd166: ff_rdata <= 8'hE1;
			14'd167: ff_rdata <= 8'hED;
			14'd168: ff_rdata <= 8'h5B;
			14'd169: ff_rdata <= 8'h80;
			14'd170: ff_rdata <= 8'h40;
			14'd171: ff_rdata <= 8'h7A;
			14'd172: ff_rdata <= 8'hA3;
			14'd173: ff_rdata <= 8'h3C;
			14'd174: ff_rdata <= 8'hD5;
			14'd175: ff_rdata <= 8'hC0;
			14'd176: ff_rdata <= 8'hD1;
			14'd177: ff_rdata <= 8'h37;
			14'd178: ff_rdata <= 8'hC9;
			14'd179: ff_rdata <= 8'h46;
			14'd180: ff_rdata <= 8'h4D;
			14'd181: ff_rdata <= 8'h50;
			14'd182: ff_rdata <= 8'h41;
			14'd183: ff_rdata <= 8'h43;
			14'd184: ff_rdata <= 8'h00;
			14'd185: ff_rdata <= 8'hFF;
			14'd186: ff_rdata <= 8'hFF;
			14'd187: ff_rdata <= 8'hFF;
			14'd188: ff_rdata <= 8'hFF;
			14'd189: ff_rdata <= 8'hFF;
			14'd190: ff_rdata <= 8'hFF;
			14'd191: ff_rdata <= 8'hFF;
			14'd192: ff_rdata <= 8'hFF;
			14'd193: ff_rdata <= 8'hFF;
			14'd194: ff_rdata <= 8'hFF;
			14'd195: ff_rdata <= 8'hFF;
			14'd196: ff_rdata <= 8'hFF;
			14'd197: ff_rdata <= 8'hFF;
			14'd198: ff_rdata <= 8'hFF;
			14'd199: ff_rdata <= 8'hFF;
			14'd200: ff_rdata <= 8'hFF;
			14'd201: ff_rdata <= 8'hFF;
			14'd202: ff_rdata <= 8'hFF;
			14'd203: ff_rdata <= 8'hFF;
			14'd204: ff_rdata <= 8'hFF;
			14'd205: ff_rdata <= 8'hFF;
			14'd206: ff_rdata <= 8'hFF;
			14'd207: ff_rdata <= 8'hFF;
			14'd208: ff_rdata <= 8'hFF;
			14'd209: ff_rdata <= 8'hFF;
			14'd210: ff_rdata <= 8'hFF;
			14'd211: ff_rdata <= 8'hFF;
			14'd212: ff_rdata <= 8'hFF;
			14'd213: ff_rdata <= 8'hFF;
			14'd214: ff_rdata <= 8'hFF;
			14'd215: ff_rdata <= 8'hFF;
			14'd216: ff_rdata <= 8'hFF;
			14'd217: ff_rdata <= 8'hFF;
			14'd218: ff_rdata <= 8'hFF;
			14'd219: ff_rdata <= 8'hFF;
			14'd220: ff_rdata <= 8'hFF;
			14'd221: ff_rdata <= 8'hFF;
			14'd222: ff_rdata <= 8'hFF;
			14'd223: ff_rdata <= 8'hFF;
			14'd224: ff_rdata <= 8'hFF;
			14'd225: ff_rdata <= 8'hFF;
			14'd226: ff_rdata <= 8'hFF;
			14'd227: ff_rdata <= 8'hFF;
			14'd228: ff_rdata <= 8'hFF;
			14'd229: ff_rdata <= 8'hFF;
			14'd230: ff_rdata <= 8'hFF;
			14'd231: ff_rdata <= 8'hFF;
			14'd232: ff_rdata <= 8'hFF;
			14'd233: ff_rdata <= 8'hFF;
			14'd234: ff_rdata <= 8'hFF;
			14'd235: ff_rdata <= 8'hFF;
			14'd236: ff_rdata <= 8'hFF;
			14'd237: ff_rdata <= 8'hFF;
			14'd238: ff_rdata <= 8'hFF;
			14'd239: ff_rdata <= 8'hFF;
			14'd240: ff_rdata <= 8'hFF;
			14'd241: ff_rdata <= 8'hFF;
			14'd242: ff_rdata <= 8'hFF;
			14'd243: ff_rdata <= 8'hFF;
			14'd244: ff_rdata <= 8'hFF;
			14'd245: ff_rdata <= 8'hFF;
			14'd246: ff_rdata <= 8'hFF;
			14'd247: ff_rdata <= 8'hFF;
			14'd248: ff_rdata <= 8'hFF;
			14'd249: ff_rdata <= 8'hFF;
			14'd250: ff_rdata <= 8'hFF;
			14'd251: ff_rdata <= 8'hFF;
			14'd252: ff_rdata <= 8'hFF;
			14'd253: ff_rdata <= 8'hFF;
			14'd254: ff_rdata <= 8'hFF;
			14'd255: ff_rdata <= 8'hFF;
			14'd256: ff_rdata <= 8'h56;
			14'd257: ff_rdata <= 8'h31;
			14'd258: ff_rdata <= 8'h2E;
			14'd259: ff_rdata <= 8'h33;
			14'd260: ff_rdata <= 8'h20;
			14'd261: ff_rdata <= 8'h31;
			14'd262: ff_rdata <= 8'h39;
			14'd263: ff_rdata <= 8'h38;
			14'd264: ff_rdata <= 8'h38;
			14'd265: ff_rdata <= 8'h20;
			14'd266: ff_rdata <= 8'h30;
			14'd267: ff_rdata <= 8'h34;
			14'd268: ff_rdata <= 8'h20;
			14'd269: ff_rdata <= 8'h32;
			14'd270: ff_rdata <= 8'h36;
			14'd271: ff_rdata <= 8'h00;
			14'd272: ff_rdata <= 8'hC3;
			14'd273: ff_rdata <= 8'h40;
			14'd274: ff_rdata <= 8'h41;
			14'd275: ff_rdata <= 8'hC3;
			14'd276: ff_rdata <= 8'h7B;
			14'd277: ff_rdata <= 8'h41;
			14'd278: ff_rdata <= 8'hC3;
			14'd279: ff_rdata <= 8'hCE;
			14'd280: ff_rdata <= 8'h42;
			14'd281: ff_rdata <= 8'hC3;
			14'd282: ff_rdata <= 8'hDA;
			14'd283: ff_rdata <= 8'h43;
			14'd284: ff_rdata <= 8'hC3;
			14'd285: ff_rdata <= 8'h30;
			14'd286: ff_rdata <= 8'h44;
			14'd287: ff_rdata <= 8'hC3;
			14'd288: ff_rdata <= 8'h47;
			14'd289: ff_rdata <= 8'h44;
			14'd290: ff_rdata <= 8'hC3;
			14'd291: ff_rdata <= 8'h3B;
			14'd292: ff_rdata <= 8'h47;
			14'd293: ff_rdata <= 8'hC9;
			14'd294: ff_rdata <= 8'h26;
			14'd295: ff_rdata <= 8'h47;
			14'd296: ff_rdata <= 8'hAB;
			14'd297: ff_rdata <= 8'h00;
			14'd298: ff_rdata <= 8'hB5;
			14'd299: ff_rdata <= 8'h00;
			14'd300: ff_rdata <= 8'hC0;
			14'd301: ff_rdata <= 8'h00;
			14'd302: ff_rdata <= 8'hCC;
			14'd303: ff_rdata <= 8'h00;
			14'd304: ff_rdata <= 8'hD8;
			14'd305: ff_rdata <= 8'h00;
			14'd306: ff_rdata <= 8'hE5;
			14'd307: ff_rdata <= 8'h00;
			14'd308: ff_rdata <= 8'hF2;
			14'd309: ff_rdata <= 8'h00;
			14'd310: ff_rdata <= 8'h01;
			14'd311: ff_rdata <= 8'h01;
			14'd312: ff_rdata <= 8'h10;
			14'd313: ff_rdata <= 8'h01;
			14'd314: ff_rdata <= 8'h20;
			14'd315: ff_rdata <= 8'h01;
			14'd316: ff_rdata <= 8'h31;
			14'd317: ff_rdata <= 8'h01;
			14'd318: ff_rdata <= 8'h43;
			14'd319: ff_rdata <= 8'h01;
			14'd320: ff_rdata <= 8'hD3;
			14'd321: ff_rdata <= 8'h7C;
			14'd322: ff_rdata <= 8'hF5;
			14'd323: ff_rdata <= 8'h7B;
			14'd324: ff_rdata <= 8'hD3;
			14'd325: ff_rdata <= 8'h7D;
			14'd326: ff_rdata <= 8'hE3;
			14'd327: ff_rdata <= 8'hE3;
			14'd328: ff_rdata <= 8'hE3;
			14'd329: ff_rdata <= 8'hE3;
			14'd330: ff_rdata <= 8'hE3;
			14'd331: ff_rdata <= 8'hE3;
			14'd332: ff_rdata <= 8'hE3;
			14'd333: ff_rdata <= 8'hE3;
			14'd334: ff_rdata <= 8'hF1;
			14'd335: ff_rdata <= 8'hC9;
			14'd336: ff_rdata <= 8'hFD;
			14'd337: ff_rdata <= 8'hE5;
			14'd338: ff_rdata <= 8'hD5;
			14'd339: ff_rdata <= 8'hC6;
			14'd340: ff_rdata <= 8'h00;
			14'd341: ff_rdata <= 8'h16;
			14'd342: ff_rdata <= 8'h00;
			14'd343: ff_rdata <= 8'h5F;
			14'd344: ff_rdata <= 8'hFD;
			14'd345: ff_rdata <= 8'h19;
			14'd346: ff_rdata <= 8'hD1;
			14'd347: ff_rdata <= 8'hD3;
			14'd348: ff_rdata <= 8'h7C;
			14'd349: ff_rdata <= 8'hF5;
			14'd350: ff_rdata <= 8'h7B;
			14'd351: ff_rdata <= 8'hD3;
			14'd352: ff_rdata <= 8'h7D;
			14'd353: ff_rdata <= 8'hFD;
			14'd354: ff_rdata <= 8'h77;
			14'd355: ff_rdata <= 8'h00;
			14'd356: ff_rdata <= 8'hE3;
			14'd357: ff_rdata <= 8'hE3;
			14'd358: ff_rdata <= 8'hE3;
			14'd359: ff_rdata <= 8'hE3;
			14'd360: ff_rdata <= 8'hF1;
			14'd361: ff_rdata <= 8'hFD;
			14'd362: ff_rdata <= 8'hE1;
			14'd363: ff_rdata <= 8'hC9;
			14'd364: ff_rdata <= 8'hE5;
			14'd365: ff_rdata <= 8'hFD;
			14'd366: ff_rdata <= 8'hE5;
			14'd367: ff_rdata <= 8'hE1;
			14'd368: ff_rdata <= 8'hC6;
			14'd369: ff_rdata <= 8'h00;
			14'd370: ff_rdata <= 8'h85;
			14'd371: ff_rdata <= 8'h6F;
			14'd372: ff_rdata <= 8'h7C;
			14'd373: ff_rdata <= 8'hCE;
			14'd374: ff_rdata <= 8'h00;
			14'd375: ff_rdata <= 8'h67;
			14'd376: ff_rdata <= 8'h7E;
			14'd377: ff_rdata <= 8'hE1;
			14'd378: ff_rdata <= 8'hC9;
			14'd379: ff_rdata <= 8'hF3;
			14'd380: ff_rdata <= 8'h7D;
			14'd381: ff_rdata <= 8'hE6;
			14'd382: ff_rdata <= 8'hFE;
			14'd383: ff_rdata <= 8'h6F;
			14'd384: ff_rdata <= 8'hE5;
			14'd385: ff_rdata <= 8'h01;
			14'd386: ff_rdata <= 8'h00;
			14'd387: ff_rdata <= 8'h40;
			14'd388: ff_rdata <= 8'hCD;
			14'd389: ff_rdata <= 8'hDC;
			14'd390: ff_rdata <= 8'h41;
			14'd391: ff_rdata <= 8'hC1;
			14'd392: ff_rdata <= 8'h7E;
			14'd393: ff_rdata <= 8'hE6;
			14'd394: ff_rdata <= 8'h01;
			14'd395: ff_rdata <= 8'hB1;
			14'd396: ff_rdata <= 8'h77;
			14'd397: ff_rdata <= 8'h23;
			14'd398: ff_rdata <= 8'h70;
			14'd399: ff_rdata <= 8'hC5;
			14'd400: ff_rdata <= 8'hFD;
			14'd401: ff_rdata <= 8'hE1;
			14'd402: ff_rdata <= 8'hCD;
			14'd403: ff_rdata <= 8'h30;
			14'd404: ff_rdata <= 8'h42;
			14'd405: ff_rdata <= 8'hFD;
			14'd406: ff_rdata <= 8'hE5;
			14'd407: ff_rdata <= 8'hE1;
			14'd408: ff_rdata <= 8'h11;
			14'd409: ff_rdata <= 8'h00;
			14'd410: ff_rdata <= 8'h00;
			14'd411: ff_rdata <= 8'h19;
			14'd412: ff_rdata <= 8'h5D;
			14'd413: ff_rdata <= 8'h54;
			14'd414: ff_rdata <= 8'h13;
			14'd415: ff_rdata <= 8'h01;
			14'd416: ff_rdata <= 8'hA0;
			14'd417: ff_rdata <= 8'h00;
			14'd418: ff_rdata <= 8'h36;
			14'd419: ff_rdata <= 8'h00;
			14'd420: ff_rdata <= 8'hED;
			14'd421: ff_rdata <= 8'hB0;
			14'd422: ff_rdata <= 8'h3E;
			14'd423: ff_rdata <= 8'h00;
			14'd424: ff_rdata <= 8'hCD;
			14'd425: ff_rdata <= 8'h3B;
			14'd426: ff_rdata <= 8'h46;
			14'd427: ff_rdata <= 8'h3E;
			14'd428: ff_rdata <= 8'h0E;
			14'd429: ff_rdata <= 8'h1E;
			14'd430: ff_rdata <= 8'h00;
			14'd431: ff_rdata <= 8'hCD;
			14'd432: ff_rdata <= 8'h50;
			14'd433: ff_rdata <= 8'h41;
			14'd434: ff_rdata <= 8'h3C;
			14'd435: ff_rdata <= 8'hCD;
			14'd436: ff_rdata <= 8'h50;
			14'd437: ff_rdata <= 8'h41;
			14'd438: ff_rdata <= 8'h3E;
			14'd439: ff_rdata <= 8'h10;
			14'd440: ff_rdata <= 8'h1E;
			14'd441: ff_rdata <= 8'h20;
			14'd442: ff_rdata <= 8'h06;
			14'd443: ff_rdata <= 8'h09;
			14'd444: ff_rdata <= 8'hCD;
			14'd445: ff_rdata <= 8'h50;
			14'd446: ff_rdata <= 8'h41;
			14'd447: ff_rdata <= 8'h3C;
			14'd448: ff_rdata <= 8'h10;
			14'd449: ff_rdata <= 8'hFA;
			14'd450: ff_rdata <= 8'h3E;
			14'd451: ff_rdata <= 8'h20;
			14'd452: ff_rdata <= 8'h1E;
			14'd453: ff_rdata <= 8'h07;
			14'd454: ff_rdata <= 8'h06;
			14'd455: ff_rdata <= 8'h09;
			14'd456: ff_rdata <= 8'hCD;
			14'd457: ff_rdata <= 8'h50;
			14'd458: ff_rdata <= 8'h41;
			14'd459: ff_rdata <= 8'h3C;
			14'd460: ff_rdata <= 8'h10;
			14'd461: ff_rdata <= 8'hFA;
			14'd462: ff_rdata <= 8'h3E;
			14'd463: ff_rdata <= 8'h30;
			14'd464: ff_rdata <= 8'h1E;
			14'd465: ff_rdata <= 8'hB3;
			14'd466: ff_rdata <= 8'h06;
			14'd467: ff_rdata <= 8'h09;
			14'd468: ff_rdata <= 8'hCD;
			14'd469: ff_rdata <= 8'h50;
			14'd470: ff_rdata <= 8'h41;
			14'd471: ff_rdata <= 8'h3C;
			14'd472: ff_rdata <= 8'h10;
			14'd473: ff_rdata <= 8'hFA;
			14'd474: ff_rdata <= 8'hFB;
			14'd475: ff_rdata <= 8'hC9;
			14'd476: ff_rdata <= 8'hCD;
			14'd477: ff_rdata <= 8'hF6;
			14'd478: ff_rdata <= 8'h41;
			14'd479: ff_rdata <= 8'hE6;
			14'd480: ff_rdata <= 8'h0F;
			14'd481: ff_rdata <= 8'h6F;
			14'd482: ff_rdata <= 8'h07;
			14'd483: ff_rdata <= 8'h07;
			14'd484: ff_rdata <= 8'h07;
			14'd485: ff_rdata <= 8'h07;
			14'd486: ff_rdata <= 8'hE6;
			14'd487: ff_rdata <= 8'h30;
			14'd488: ff_rdata <= 8'hB5;
			14'd489: ff_rdata <= 8'hE6;
			14'd490: ff_rdata <= 8'h3C;
			14'd491: ff_rdata <= 8'hF6;
			14'd492: ff_rdata <= 8'h01;
			14'd493: ff_rdata <= 8'h07;
			14'd494: ff_rdata <= 8'h5F;
			14'd495: ff_rdata <= 8'h16;
			14'd496: ff_rdata <= 8'h00;
			14'd497: ff_rdata <= 8'h21;
			14'd498: ff_rdata <= 8'h09;
			14'd499: ff_rdata <= 8'hFD;
			14'd500: ff_rdata <= 8'h19;
			14'd501: ff_rdata <= 8'hC9;
			14'd502: ff_rdata <= 8'hC5;
			14'd503: ff_rdata <= 8'hD5;
			14'd504: ff_rdata <= 8'hE5;
			14'd505: ff_rdata <= 8'h78;
			14'd506: ff_rdata <= 8'h07;
			14'd507: ff_rdata <= 8'h07;
			14'd508: ff_rdata <= 8'hE6;
			14'd509: ff_rdata <= 8'h03;
			14'd510: ff_rdata <= 8'h47;
			14'd511: ff_rdata <= 8'hDB;
			14'd512: ff_rdata <= 8'hA8;
			14'd513: ff_rdata <= 8'hCD;
			14'd514: ff_rdata <= 8'h26;
			14'd515: ff_rdata <= 8'h42;
			14'd516: ff_rdata <= 8'hE6;
			14'd517: ff_rdata <= 8'h03;
			14'd518: ff_rdata <= 8'h5F;
			14'd519: ff_rdata <= 8'h16;
			14'd520: ff_rdata <= 8'h00;
			14'd521: ff_rdata <= 8'h21;
			14'd522: ff_rdata <= 8'hC1;
			14'd523: ff_rdata <= 8'hFC;
			14'd524: ff_rdata <= 8'h19;
			14'd525: ff_rdata <= 8'h7E;
			14'd526: ff_rdata <= 8'hE6;
			14'd527: ff_rdata <= 8'h80;
			14'd528: ff_rdata <= 8'hB3;
			14'd529: ff_rdata <= 8'hF2;
			14'd530: ff_rdata <= 8'h22;
			14'd531: ff_rdata <= 8'h42;
			14'd532: ff_rdata <= 8'h5F;
			14'd533: ff_rdata <= 8'h23;
			14'd534: ff_rdata <= 8'h23;
			14'd535: ff_rdata <= 8'h23;
			14'd536: ff_rdata <= 8'h23;
			14'd537: ff_rdata <= 8'h7E;
			14'd538: ff_rdata <= 8'h07;
			14'd539: ff_rdata <= 8'h07;
			14'd540: ff_rdata <= 8'hCD;
			14'd541: ff_rdata <= 8'h26;
			14'd542: ff_rdata <= 8'h42;
			14'd543: ff_rdata <= 8'hE6;
			14'd544: ff_rdata <= 8'h0C;
			14'd545: ff_rdata <= 8'hB3;
			14'd546: ff_rdata <= 8'hE1;
			14'd547: ff_rdata <= 8'hD1;
			14'd548: ff_rdata <= 8'hC1;
			14'd549: ff_rdata <= 8'hC9;
			14'd550: ff_rdata <= 8'h04;
			14'd551: ff_rdata <= 8'h05;
			14'd552: ff_rdata <= 8'hC8;
			14'd553: ff_rdata <= 8'hC5;
			14'd554: ff_rdata <= 8'h0F;
			14'd555: ff_rdata <= 8'h0F;
			14'd556: ff_rdata <= 8'h10;
			14'd557: ff_rdata <= 8'hFC;
			14'd558: ff_rdata <= 8'hC1;
			14'd559: ff_rdata <= 8'hC9;
			14'd560: ff_rdata <= 8'h21;
			14'd561: ff_rdata <= 8'h43;
			14'd562: ff_rdata <= 8'h42;
			14'd563: ff_rdata <= 8'hFD;
			14'd564: ff_rdata <= 8'hE5;
			14'd565: ff_rdata <= 8'hD1;
			14'd566: ff_rdata <= 8'h01;
			14'd567: ff_rdata <= 8'h8B;
			14'd568: ff_rdata <= 8'h00;
			14'd569: ff_rdata <= 8'hED;
			14'd570: ff_rdata <= 8'hB0;
			14'd571: ff_rdata <= 8'h01;
			14'd572: ff_rdata <= 8'h00;
			14'd573: ff_rdata <= 8'h40;
			14'd574: ff_rdata <= 8'hCD;
			14'd575: ff_rdata <= 8'hF6;
			14'd576: ff_rdata <= 8'h41;
			14'd577: ff_rdata <= 8'hFD;
			14'd578: ff_rdata <= 8'hE9;
			14'd579: ff_rdata <= 8'hF5;
			14'd580: ff_rdata <= 8'hFD;
			14'd581: ff_rdata <= 8'hE5;
			14'd582: ff_rdata <= 8'hD1;
			14'd583: ff_rdata <= 8'h21;
			14'd584: ff_rdata <= 8'h15;
			14'd585: ff_rdata <= 8'h00;
			14'd586: ff_rdata <= 8'h19;
			14'd587: ff_rdata <= 8'hE5;
			14'd588: ff_rdata <= 8'h21;
			14'd589: ff_rdata <= 8'h7B;
			14'd590: ff_rdata <= 8'h00;
			14'd591: ff_rdata <= 8'h19;
			14'd592: ff_rdata <= 8'hDD;
			14'd593: ff_rdata <= 8'h21;
			14'd594: ff_rdata <= 8'h37;
			14'd595: ff_rdata <= 8'h00;
			14'd596: ff_rdata <= 8'hDD;
			14'd597: ff_rdata <= 8'h19;
			14'd598: ff_rdata <= 8'hDD;
			14'd599: ff_rdata <= 8'hE9;
			14'd600: ff_rdata <= 8'hFE;
			14'd601: ff_rdata <= 8'hFF;
			14'd602: ff_rdata <= 8'h20;
			14'd603: ff_rdata <= 8'h16;
			14'd604: ff_rdata <= 8'hFD;
			14'd605: ff_rdata <= 8'hE5;
			14'd606: ff_rdata <= 8'hD1;
			14'd607: ff_rdata <= 8'h21;
			14'd608: ff_rdata <= 8'h27;
			14'd609: ff_rdata <= 8'h00;
			14'd610: ff_rdata <= 8'h19;
			14'd611: ff_rdata <= 8'hE5;
			14'd612: ff_rdata <= 8'h21;
			14'd613: ff_rdata <= 8'h83;
			14'd614: ff_rdata <= 8'h00;
			14'd615: ff_rdata <= 8'h19;
			14'd616: ff_rdata <= 8'hDD;
			14'd617: ff_rdata <= 8'hE9;
			14'd618: ff_rdata <= 8'h3A;
			14'd619: ff_rdata <= 8'hF6;
			14'd620: ff_rdata <= 8'h7F;
			14'd621: ff_rdata <= 8'hF6;
			14'd622: ff_rdata <= 8'h01;
			14'd623: ff_rdata <= 8'h32;
			14'd624: ff_rdata <= 8'hF6;
			14'd625: ff_rdata <= 8'h7F;
			14'd626: ff_rdata <= 8'hF1;
			14'd627: ff_rdata <= 8'h21;
			14'd628: ff_rdata <= 8'h00;
			14'd629: ff_rdata <= 8'h40;
			14'd630: ff_rdata <= 8'hCD;
			14'd631: ff_rdata <= 8'h24;
			14'd632: ff_rdata <= 8'h00;
			14'd633: ff_rdata <= 8'hC9;
			14'd634: ff_rdata <= 8'hEB;
			14'd635: ff_rdata <= 8'h21;
			14'd636: ff_rdata <= 8'hC1;
			14'd637: ff_rdata <= 8'hFC;
			14'd638: ff_rdata <= 8'h0E;
			14'd639: ff_rdata <= 8'h00;
			14'd640: ff_rdata <= 8'h06;
			14'd641: ff_rdata <= 8'h04;
			14'd642: ff_rdata <= 8'hC5;
			14'd643: ff_rdata <= 8'hE5;
			14'd644: ff_rdata <= 8'h7E;
			14'd645: ff_rdata <= 8'hE6;
			14'd646: ff_rdata <= 8'h80;
			14'd647: ff_rdata <= 8'hB1;
			14'd648: ff_rdata <= 8'h4F;
			14'd649: ff_rdata <= 8'h06;
			14'd650: ff_rdata <= 8'h01;
			14'd651: ff_rdata <= 8'h07;
			14'd652: ff_rdata <= 8'h30;
			14'd653: ff_rdata <= 8'h02;
			14'd654: ff_rdata <= 8'h06;
			14'd655: ff_rdata <= 8'h04;
			14'd656: ff_rdata <= 8'hC5;
			14'd657: ff_rdata <= 8'hD5;
			14'd658: ff_rdata <= 8'h79;
			14'd659: ff_rdata <= 8'h26;
			14'd660: ff_rdata <= 8'h40;
			14'd661: ff_rdata <= 8'hCD;
			14'd662: ff_rdata <= 8'h24;
			14'd663: ff_rdata <= 8'h00;
			14'd664: ff_rdata <= 8'hD1;
			14'd665: ff_rdata <= 8'hD5;
			14'd666: ff_rdata <= 8'h21;
			14'd667: ff_rdata <= 8'h18;
			14'd668: ff_rdata <= 8'h40;
			14'd669: ff_rdata <= 8'h06;
			14'd670: ff_rdata <= 8'h08;
			14'd671: ff_rdata <= 8'h1A;
			14'd672: ff_rdata <= 8'h13;
			14'd673: ff_rdata <= 8'hBE;
			14'd674: ff_rdata <= 8'h23;
			14'd675: ff_rdata <= 8'h20;
			14'd676: ff_rdata <= 8'h02;
			14'd677: ff_rdata <= 8'h10;
			14'd678: ff_rdata <= 8'hF8;
			14'd679: ff_rdata <= 8'hD1;
			14'd680: ff_rdata <= 8'hC1;
			14'd681: ff_rdata <= 8'h28;
			14'd682: ff_rdata <= 8'h0F;
			14'd683: ff_rdata <= 8'h79;
			14'd684: ff_rdata <= 8'hC6;
			14'd685: ff_rdata <= 8'h04;
			14'd686: ff_rdata <= 8'h4F;
			14'd687: ff_rdata <= 8'h10;
			14'd688: ff_rdata <= 8'hDF;
			14'd689: ff_rdata <= 8'hE1;
			14'd690: ff_rdata <= 8'hC1;
			14'd691: ff_rdata <= 8'h23;
			14'd692: ff_rdata <= 8'h0C;
			14'd693: ff_rdata <= 8'h10;
			14'd694: ff_rdata <= 8'hCB;
			14'd695: ff_rdata <= 8'h3E;
			14'd696: ff_rdata <= 8'hFF;
			14'd697: ff_rdata <= 8'hC9;
			14'd698: ff_rdata <= 8'h79;
			14'd699: ff_rdata <= 8'hE1;
			14'd700: ff_rdata <= 8'hC1;
			14'd701: ff_rdata <= 8'hC9;
			14'd702: ff_rdata <= 8'h41;
			14'd703: ff_rdata <= 8'h50;
			14'd704: ff_rdata <= 8'h52;
			14'd705: ff_rdata <= 8'h4C;
			14'd706: ff_rdata <= 8'h4F;
			14'd707: ff_rdata <= 8'h50;
			14'd708: ff_rdata <= 8'h4C;
			14'd709: ff_rdata <= 8'h4C;
			14'd710: ff_rdata <= 8'h50;
			14'd711: ff_rdata <= 8'h41;
			14'd712: ff_rdata <= 8'h43;
			14'd713: ff_rdata <= 8'h32;
			14'd714: ff_rdata <= 8'h4F;
			14'd715: ff_rdata <= 8'h50;
			14'd716: ff_rdata <= 8'h4C;
			14'd717: ff_rdata <= 8'h4C;
			14'd718: ff_rdata <= 8'hF3;
			14'd719: ff_rdata <= 8'hE5;
			14'd720: ff_rdata <= 8'hF5;
			14'd721: ff_rdata <= 8'h01;
			14'd722: ff_rdata <= 8'h00;
			14'd723: ff_rdata <= 8'h40;
			14'd724: ff_rdata <= 8'hCD;
			14'd725: ff_rdata <= 8'hDC;
			14'd726: ff_rdata <= 8'h41;
			14'd727: ff_rdata <= 8'h7E;
			14'd728: ff_rdata <= 8'h23;
			14'd729: ff_rdata <= 8'h66;
			14'd730: ff_rdata <= 8'hE6;
			14'd731: ff_rdata <= 8'hFE;
			14'd732: ff_rdata <= 8'h6F;
			14'd733: ff_rdata <= 8'hE5;
			14'd734: ff_rdata <= 8'hFD;
			14'd735: ff_rdata <= 8'hE1;
			14'd736: ff_rdata <= 8'h11;
			14'd737: ff_rdata <= 8'h3D;
			14'd738: ff_rdata <= 8'h00;
			14'd739: ff_rdata <= 8'h19;
			14'd740: ff_rdata <= 8'hE5;
			14'd741: ff_rdata <= 8'hDD;
			14'd742: ff_rdata <= 8'hE1;
			14'd743: ff_rdata <= 8'hF1;
			14'd744: ff_rdata <= 8'hB7;
			14'd745: ff_rdata <= 8'h20;
			14'd746: ff_rdata <= 8'h01;
			14'd747: ff_rdata <= 8'h3D;
			14'd748: ff_rdata <= 8'hFD;
			14'd749: ff_rdata <= 8'h77;
			14'd750: ff_rdata <= 8'h3A;
			14'd751: ff_rdata <= 8'hE1;
			14'd752: ff_rdata <= 8'h7E;
			14'd753: ff_rdata <= 8'hFE;
			14'd754: ff_rdata <= 8'h12;
			14'd755: ff_rdata <= 8'hC2;
			14'd756: ff_rdata <= 8'h06;
			14'd757: ff_rdata <= 8'h43;
			14'd758: ff_rdata <= 8'h3E;
			14'd759: ff_rdata <= 8'h0E;
			14'd760: ff_rdata <= 8'h1E;
			14'd761: ff_rdata <= 8'h00;
			14'd762: ff_rdata <= 8'hCD;
			14'd763: ff_rdata <= 8'h50;
			14'd764: ff_rdata <= 8'h41;
			14'd765: ff_rdata <= 8'h06;
			14'd766: ff_rdata <= 8'h09;
			14'd767: ff_rdata <= 8'hFD;
			14'd768: ff_rdata <= 8'h36;
			14'd769: ff_rdata <= 8'h39;
			14'd770: ff_rdata <= 8'h00;
			14'd771: ff_rdata <= 8'hC3;
			14'd772: ff_rdata <= 8'h0C;
			14'd773: ff_rdata <= 8'h43;
			14'd774: ff_rdata <= 8'h06;
			14'd775: ff_rdata <= 8'h07;
			14'd776: ff_rdata <= 8'hFD;
			14'd777: ff_rdata <= 8'h36;
			14'd778: ff_rdata <= 8'h39;
			14'd779: ff_rdata <= 8'hFF;
			14'd780: ff_rdata <= 8'hFD;
			14'd781: ff_rdata <= 8'h36;
			14'd782: ff_rdata <= 8'h3B;
			14'd783: ff_rdata <= 8'h00;
			14'd784: ff_rdata <= 8'hE5;
			14'd785: ff_rdata <= 8'h5E;
			14'd786: ff_rdata <= 8'h23;
			14'd787: ff_rdata <= 8'h56;
			14'd788: ff_rdata <= 8'h23;
			14'd789: ff_rdata <= 8'h7A;
			14'd790: ff_rdata <= 8'hB3;
			14'd791: ff_rdata <= 8'hC2;
			14'd792: ff_rdata <= 8'h25;
			14'd793: ff_rdata <= 8'h43;
			14'd794: ff_rdata <= 8'hDD;
			14'd795: ff_rdata <= 8'h36;
			14'd796: ff_rdata <= 8'h00;
			14'd797: ff_rdata <= 8'h00;
			14'd798: ff_rdata <= 8'hDD;
			14'd799: ff_rdata <= 8'h36;
			14'd800: ff_rdata <= 8'h01;
			14'd801: ff_rdata <= 8'h00;
			14'd802: ff_rdata <= 8'hC3;
			14'd803: ff_rdata <= 8'h37;
			14'd804: ff_rdata <= 8'h43;
			14'd805: ff_rdata <= 8'hE3;
			14'd806: ff_rdata <= 8'hEB;
			14'd807: ff_rdata <= 8'h19;
			14'd808: ff_rdata <= 8'hDD;
			14'd809: ff_rdata <= 8'h75;
			14'd810: ff_rdata <= 8'h00;
			14'd811: ff_rdata <= 8'hDD;
			14'd812: ff_rdata <= 8'h74;
			14'd813: ff_rdata <= 8'h01;
			14'd814: ff_rdata <= 8'hDD;
			14'd815: ff_rdata <= 8'h36;
			14'd816: ff_rdata <= 8'h0A;
			14'd817: ff_rdata <= 8'h01;
			14'd818: ff_rdata <= 8'hEB;
			14'd819: ff_rdata <= 8'hE3;
			14'd820: ff_rdata <= 8'hFD;
			14'd821: ff_rdata <= 8'h34;
			14'd822: ff_rdata <= 8'h3B;
			14'd823: ff_rdata <= 8'h11;
			14'd824: ff_rdata <= 8'h0B;
			14'd825: ff_rdata <= 8'h00;
			14'd826: ff_rdata <= 8'hDD;
			14'd827: ff_rdata <= 8'h19;
			14'd828: ff_rdata <= 8'h10;
			14'd829: ff_rdata <= 8'hD3;
			14'd830: ff_rdata <= 8'hE1;
			14'd831: ff_rdata <= 8'hCD;
			14'd832: ff_rdata <= 8'h44;
			14'd833: ff_rdata <= 8'h43;
			14'd834: ff_rdata <= 8'hFB;
			14'd835: ff_rdata <= 8'hC9;
			14'd836: ff_rdata <= 8'hFD;
			14'd837: ff_rdata <= 8'hE5;
			14'd838: ff_rdata <= 8'hDD;
			14'd839: ff_rdata <= 8'hE1;
			14'd840: ff_rdata <= 8'h11;
			14'd841: ff_rdata <= 8'h3D;
			14'd842: ff_rdata <= 8'h00;
			14'd843: ff_rdata <= 8'hDD;
			14'd844: ff_rdata <= 8'h19;
			14'd845: ff_rdata <= 8'h06;
			14'd846: ff_rdata <= 8'h09;
			14'd847: ff_rdata <= 8'hFD;
			14'd848: ff_rdata <= 8'h7E;
			14'd849: ff_rdata <= 8'h39;
			14'd850: ff_rdata <= 8'hB7;
			14'd851: ff_rdata <= 8'hCA;
			14'd852: ff_rdata <= 8'h74;
			14'd853: ff_rdata <= 8'h43;
			14'd854: ff_rdata <= 8'hDD;
			14'd855: ff_rdata <= 8'h6E;
			14'd856: ff_rdata <= 8'h00;
			14'd857: ff_rdata <= 8'hDD;
			14'd858: ff_rdata <= 8'h66;
			14'd859: ff_rdata <= 8'h01;
			14'd860: ff_rdata <= 8'hDD;
			14'd861: ff_rdata <= 8'h75;
			14'd862: ff_rdata <= 8'h02;
			14'd863: ff_rdata <= 8'hDD;
			14'd864: ff_rdata <= 8'h74;
			14'd865: ff_rdata <= 8'h03;
			14'd866: ff_rdata <= 8'hDD;
			14'd867: ff_rdata <= 8'h36;
			14'd868: ff_rdata <= 8'h04;
			14'd869: ff_rdata <= 8'h01;
			14'd870: ff_rdata <= 8'hDD;
			14'd871: ff_rdata <= 8'h36;
			14'd872: ff_rdata <= 8'h05;
			14'd873: ff_rdata <= 8'h00;
			14'd874: ff_rdata <= 8'hCD;
			14'd875: ff_rdata <= 8'hB5;
			14'd876: ff_rdata <= 8'h43;
			14'd877: ff_rdata <= 8'h11;
			14'd878: ff_rdata <= 8'h0B;
			14'd879: ff_rdata <= 8'h00;
			14'd880: ff_rdata <= 8'hDD;
			14'd881: ff_rdata <= 8'h19;
			14'd882: ff_rdata <= 8'h06;
			14'd883: ff_rdata <= 8'h06;
			14'd884: ff_rdata <= 8'hDD;
			14'd885: ff_rdata <= 8'h6E;
			14'd886: ff_rdata <= 8'h00;
			14'd887: ff_rdata <= 8'hDD;
			14'd888: ff_rdata <= 8'h66;
			14'd889: ff_rdata <= 8'h01;
			14'd890: ff_rdata <= 8'hDD;
			14'd891: ff_rdata <= 8'h75;
			14'd892: ff_rdata <= 8'h02;
			14'd893: ff_rdata <= 8'hDD;
			14'd894: ff_rdata <= 8'h74;
			14'd895: ff_rdata <= 8'h03;
			14'd896: ff_rdata <= 8'hDD;
			14'd897: ff_rdata <= 8'h36;
			14'd898: ff_rdata <= 8'h04;
			14'd899: ff_rdata <= 8'h01;
			14'd900: ff_rdata <= 8'hDD;
			14'd901: ff_rdata <= 8'h36;
			14'd902: ff_rdata <= 8'h05;
			14'd903: ff_rdata <= 8'h00;
			14'd904: ff_rdata <= 8'hDD;
			14'd905: ff_rdata <= 8'h36;
			14'd906: ff_rdata <= 8'h06;
			14'd907: ff_rdata <= 8'h00;
			14'd908: ff_rdata <= 8'hDD;
			14'd909: ff_rdata <= 8'h36;
			14'd910: ff_rdata <= 8'h07;
			14'd911: ff_rdata <= 8'h00;
			14'd912: ff_rdata <= 8'hDD;
			14'd913: ff_rdata <= 8'h36;
			14'd914: ff_rdata <= 8'h09;
			14'd915: ff_rdata <= 8'h00;
			14'd916: ff_rdata <= 8'hDD;
			14'd917: ff_rdata <= 8'h36;
			14'd918: ff_rdata <= 8'h08;
			14'd919: ff_rdata <= 8'h08;
			14'd920: ff_rdata <= 8'h3E;
			14'd921: ff_rdata <= 8'h1F;
			14'd922: ff_rdata <= 8'h80;
			14'd923: ff_rdata <= 8'hCD;
			14'd924: ff_rdata <= 8'h6C;
			14'd925: ff_rdata <= 8'h41;
			14'd926: ff_rdata <= 8'hE6;
			14'd927: ff_rdata <= 8'hCF;
			14'd928: ff_rdata <= 8'h5F;
			14'd929: ff_rdata <= 8'h3E;
			14'd930: ff_rdata <= 8'h1F;
			14'd931: ff_rdata <= 8'h80;
			14'd932: ff_rdata <= 8'hCD;
			14'd933: ff_rdata <= 8'h50;
			14'd934: ff_rdata <= 8'h41;
			14'd935: ff_rdata <= 8'h11;
			14'd936: ff_rdata <= 8'h0B;
			14'd937: ff_rdata <= 8'h00;
			14'd938: ff_rdata <= 8'hDD;
			14'd939: ff_rdata <= 8'h19;
			14'd940: ff_rdata <= 8'h10;
			14'd941: ff_rdata <= 8'hC6;
			14'd942: ff_rdata <= 8'hFD;
			14'd943: ff_rdata <= 8'h7E;
			14'd944: ff_rdata <= 8'h3B;
			14'd945: ff_rdata <= 8'hFD;
			14'd946: ff_rdata <= 8'h77;
			14'd947: ff_rdata <= 8'h3C;
			14'd948: ff_rdata <= 8'hC9;
			14'd949: ff_rdata <= 8'h21;
			14'd950: ff_rdata <= 8'hC5;
			14'd951: ff_rdata <= 8'h43;
			14'd952: ff_rdata <= 8'h7E;
			14'd953: ff_rdata <= 8'hFE;
			14'd954: ff_rdata <= 8'hFF;
			14'd955: ff_rdata <= 8'hC8;
			14'd956: ff_rdata <= 8'h23;
			14'd957: ff_rdata <= 8'h5E;
			14'd958: ff_rdata <= 8'h23;
			14'd959: ff_rdata <= 8'hCD;
			14'd960: ff_rdata <= 8'h50;
			14'd961: ff_rdata <= 8'h41;
			14'd962: ff_rdata <= 8'hC3;
			14'd963: ff_rdata <= 8'hB8;
			14'd964: ff_rdata <= 8'h43;
			14'd965: ff_rdata <= 8'h0E;
			14'd966: ff_rdata <= 8'h20;
			14'd967: ff_rdata <= 8'h16;
			14'd968: ff_rdata <= 8'h20;
			14'd969: ff_rdata <= 8'h17;
			14'd970: ff_rdata <= 8'h50;
			14'd971: ff_rdata <= 8'h18;
			14'd972: ff_rdata <= 8'hC0;
			14'd973: ff_rdata <= 8'h26;
			14'd974: ff_rdata <= 8'h05;
			14'd975: ff_rdata <= 8'h27;
			14'd976: ff_rdata <= 8'h05;
			14'd977: ff_rdata <= 8'h28;
			14'd978: ff_rdata <= 8'h01;
			14'd979: ff_rdata <= 8'h36;
			14'd980: ff_rdata <= 8'h03;
			14'd981: ff_rdata <= 8'h37;
			14'd982: ff_rdata <= 8'h33;
			14'd983: ff_rdata <= 8'h38;
			14'd984: ff_rdata <= 8'h33;
			14'd985: ff_rdata <= 8'hFF;
			14'd986: ff_rdata <= 8'hF3;
			14'd987: ff_rdata <= 8'h01;
			14'd988: ff_rdata <= 8'h00;
			14'd989: ff_rdata <= 8'h40;
			14'd990: ff_rdata <= 8'hCD;
			14'd991: ff_rdata <= 8'hDC;
			14'd992: ff_rdata <= 8'h41;
			14'd993: ff_rdata <= 8'h7E;
			14'd994: ff_rdata <= 8'h23;
			14'd995: ff_rdata <= 8'h66;
			14'd996: ff_rdata <= 8'hE6;
			14'd997: ff_rdata <= 8'hFE;
			14'd998: ff_rdata <= 8'h6F;
			14'd999: ff_rdata <= 8'hE5;
			14'd1000: ff_rdata <= 8'hFD;
			14'd1001: ff_rdata <= 8'hE1;
			14'd1002: ff_rdata <= 8'h11;
			14'd1003: ff_rdata <= 8'h3D;
			14'd1004: ff_rdata <= 8'h00;
			14'd1005: ff_rdata <= 8'h19;
			14'd1006: ff_rdata <= 8'hE5;
			14'd1007: ff_rdata <= 8'hDD;
			14'd1008: ff_rdata <= 8'hE1;
			14'd1009: ff_rdata <= 8'h06;
			14'd1010: ff_rdata <= 8'h09;
			14'd1011: ff_rdata <= 8'hFD;
			14'd1012: ff_rdata <= 8'h7E;
			14'd1013: ff_rdata <= 8'h39;
			14'd1014: ff_rdata <= 8'hB7;
			14'd1015: ff_rdata <= 8'hCA;
			14'd1016: ff_rdata <= 8'h10;
			14'd1017: ff_rdata <= 8'h44;
			14'd1018: ff_rdata <= 8'h3E;
			14'd1019: ff_rdata <= 8'h0E;
			14'd1020: ff_rdata <= 8'h1E;
			14'd1021: ff_rdata <= 8'h20;
			14'd1022: ff_rdata <= 8'hCD;
			14'd1023: ff_rdata <= 8'h50;
			14'd1024: ff_rdata <= 8'h41;
			14'd1025: ff_rdata <= 8'hDD;
			14'd1026: ff_rdata <= 8'h36;
			14'd1027: ff_rdata <= 8'h02;
			14'd1028: ff_rdata <= 8'h00;
			14'd1029: ff_rdata <= 8'hDD;
			14'd1030: ff_rdata <= 8'h36;
			14'd1031: ff_rdata <= 8'h03;
			14'd1032: ff_rdata <= 8'h00;
			14'd1033: ff_rdata <= 8'h11;
			14'd1034: ff_rdata <= 8'h0B;
			14'd1035: ff_rdata <= 8'h00;
			14'd1036: ff_rdata <= 8'hDD;
			14'd1037: ff_rdata <= 8'h19;
			14'd1038: ff_rdata <= 8'h06;
			14'd1039: ff_rdata <= 8'h06;
			14'd1040: ff_rdata <= 8'hDD;
			14'd1041: ff_rdata <= 8'h36;
			14'd1042: ff_rdata <= 8'h02;
			14'd1043: ff_rdata <= 8'h00;
			14'd1044: ff_rdata <= 8'hDD;
			14'd1045: ff_rdata <= 8'h36;
			14'd1046: ff_rdata <= 8'h03;
			14'd1047: ff_rdata <= 8'h00;
			14'd1048: ff_rdata <= 8'h3E;
			14'd1049: ff_rdata <= 8'h1F;
			14'd1050: ff_rdata <= 8'h80;
			14'd1051: ff_rdata <= 8'hCD;
			14'd1052: ff_rdata <= 8'h6C;
			14'd1053: ff_rdata <= 8'h41;
			14'd1054: ff_rdata <= 8'hE6;
			14'd1055: ff_rdata <= 8'hEF;
			14'd1056: ff_rdata <= 8'h5F;
			14'd1057: ff_rdata <= 8'h3E;
			14'd1058: ff_rdata <= 8'h1F;
			14'd1059: ff_rdata <= 8'h80;
			14'd1060: ff_rdata <= 8'hCD;
			14'd1061: ff_rdata <= 8'h50;
			14'd1062: ff_rdata <= 8'h41;
			14'd1063: ff_rdata <= 8'h11;
			14'd1064: ff_rdata <= 8'h0B;
			14'd1065: ff_rdata <= 8'h00;
			14'd1066: ff_rdata <= 8'hDD;
			14'd1067: ff_rdata <= 8'h19;
			14'd1068: ff_rdata <= 8'h10;
			14'd1069: ff_rdata <= 8'hE2;
			14'd1070: ff_rdata <= 8'hFB;
			14'd1071: ff_rdata <= 8'hC9;
			14'd1072: ff_rdata <= 8'hC5;
			14'd1073: ff_rdata <= 8'hD5;
			14'd1074: ff_rdata <= 8'hE5;
			14'd1075: ff_rdata <= 8'hEB;
			14'd1076: ff_rdata <= 8'h6F;
			14'd1077: ff_rdata <= 8'h26;
			14'd1078: ff_rdata <= 8'h00;
			14'd1079: ff_rdata <= 8'h29;
			14'd1080: ff_rdata <= 8'h29;
			14'd1081: ff_rdata <= 8'h29;
			14'd1082: ff_rdata <= 8'h01;
			14'd1083: ff_rdata <= 8'h00;
			14'd1084: ff_rdata <= 8'h4C;
			14'd1085: ff_rdata <= 8'h09;
			14'd1086: ff_rdata <= 8'h01;
			14'd1087: ff_rdata <= 8'h08;
			14'd1088: ff_rdata <= 8'h00;
			14'd1089: ff_rdata <= 8'hED;
			14'd1090: ff_rdata <= 8'hB0;
			14'd1091: ff_rdata <= 8'hE1;
			14'd1092: ff_rdata <= 8'hD1;
			14'd1093: ff_rdata <= 8'hC1;
			14'd1094: ff_rdata <= 8'hC9;
			14'd1095: ff_rdata <= 8'hF5;
			14'd1096: ff_rdata <= 8'hC5;
			14'd1097: ff_rdata <= 8'hD5;
			14'd1098: ff_rdata <= 8'hE5;
			14'd1099: ff_rdata <= 8'hDD;
			14'd1100: ff_rdata <= 8'hE5;
			14'd1101: ff_rdata <= 8'hFD;
			14'd1102: ff_rdata <= 8'hE5;
			14'd1103: ff_rdata <= 8'h01;
			14'd1104: ff_rdata <= 8'h00;
			14'd1105: ff_rdata <= 8'h40;
			14'd1106: ff_rdata <= 8'hCD;
			14'd1107: ff_rdata <= 8'hDC;
			14'd1108: ff_rdata <= 8'h41;
			14'd1109: ff_rdata <= 8'h7E;
			14'd1110: ff_rdata <= 8'h23;
			14'd1111: ff_rdata <= 8'h66;
			14'd1112: ff_rdata <= 8'hE6;
			14'd1113: ff_rdata <= 8'hFE;
			14'd1114: ff_rdata <= 8'h6F;
			14'd1115: ff_rdata <= 8'hE5;
			14'd1116: ff_rdata <= 8'hFD;
			14'd1117: ff_rdata <= 8'hE1;
			14'd1118: ff_rdata <= 8'h11;
			14'd1119: ff_rdata <= 8'h3D;
			14'd1120: ff_rdata <= 8'h00;
			14'd1121: ff_rdata <= 8'h19;
			14'd1122: ff_rdata <= 8'hE5;
			14'd1123: ff_rdata <= 8'hDD;
			14'd1124: ff_rdata <= 8'hE1;
			14'd1125: ff_rdata <= 8'h06;
			14'd1126: ff_rdata <= 8'h09;
			14'd1127: ff_rdata <= 8'hFD;
			14'd1128: ff_rdata <= 8'h7E;
			14'd1129: ff_rdata <= 8'h39;
			14'd1130: ff_rdata <= 8'hB7;
			14'd1131: ff_rdata <= 8'hCA;
			14'd1132: ff_rdata <= 8'h92;
			14'd1133: ff_rdata <= 8'h44;
			14'd1134: ff_rdata <= 8'hDD;
			14'd1135: ff_rdata <= 8'h6E;
			14'd1136: ff_rdata <= 8'h02;
			14'd1137: ff_rdata <= 8'hDD;
			14'd1138: ff_rdata <= 8'h66;
			14'd1139: ff_rdata <= 8'h03;
			14'd1140: ff_rdata <= 8'h7D;
			14'd1141: ff_rdata <= 8'hB4;
			14'd1142: ff_rdata <= 8'hCA;
			14'd1143: ff_rdata <= 8'h8B;
			14'd1144: ff_rdata <= 8'h44;
			14'd1145: ff_rdata <= 8'hDD;
			14'd1146: ff_rdata <= 8'h5E;
			14'd1147: ff_rdata <= 8'h04;
			14'd1148: ff_rdata <= 8'hDD;
			14'd1149: ff_rdata <= 8'h56;
			14'd1150: ff_rdata <= 8'h05;
			14'd1151: ff_rdata <= 8'h1B;
			14'd1152: ff_rdata <= 8'h7B;
			14'd1153: ff_rdata <= 8'hB2;
			14'd1154: ff_rdata <= 8'hCC;
			14'd1155: ff_rdata <= 8'h81;
			14'd1156: ff_rdata <= 8'h46;
			14'd1157: ff_rdata <= 8'hDD;
			14'd1158: ff_rdata <= 8'h73;
			14'd1159: ff_rdata <= 8'h04;
			14'd1160: ff_rdata <= 8'hDD;
			14'd1161: ff_rdata <= 8'h72;
			14'd1162: ff_rdata <= 8'h05;
			14'd1163: ff_rdata <= 8'h11;
			14'd1164: ff_rdata <= 8'h0B;
			14'd1165: ff_rdata <= 8'h00;
			14'd1166: ff_rdata <= 8'hDD;
			14'd1167: ff_rdata <= 8'h19;
			14'd1168: ff_rdata <= 8'h06;
			14'd1169: ff_rdata <= 8'h06;
			14'd1170: ff_rdata <= 8'hDD;
			14'd1171: ff_rdata <= 8'h5E;
			14'd1172: ff_rdata <= 8'h06;
			14'd1173: ff_rdata <= 8'hDD;
			14'd1174: ff_rdata <= 8'h56;
			14'd1175: ff_rdata <= 8'h07;
			14'd1176: ff_rdata <= 8'h7B;
			14'd1177: ff_rdata <= 8'hB2;
			14'd1178: ff_rdata <= 8'hCA;
			14'd1179: ff_rdata <= 8'hA9;
			14'd1180: ff_rdata <= 8'h44;
			14'd1181: ff_rdata <= 8'h1B;
			14'd1182: ff_rdata <= 8'h7B;
			14'd1183: ff_rdata <= 8'hB2;
			14'd1184: ff_rdata <= 8'hDD;
			14'd1185: ff_rdata <= 8'h73;
			14'd1186: ff_rdata <= 8'h06;
			14'd1187: ff_rdata <= 8'hDD;
			14'd1188: ff_rdata <= 8'h72;
			14'd1189: ff_rdata <= 8'h07;
			14'd1190: ff_rdata <= 8'hCC;
			14'd1191: ff_rdata <= 8'hD6;
			14'd1192: ff_rdata <= 8'h44;
			14'd1193: ff_rdata <= 8'hDD;
			14'd1194: ff_rdata <= 8'h6E;
			14'd1195: ff_rdata <= 8'h02;
			14'd1196: ff_rdata <= 8'hDD;
			14'd1197: ff_rdata <= 8'h66;
			14'd1198: ff_rdata <= 8'h03;
			14'd1199: ff_rdata <= 8'h7D;
			14'd1200: ff_rdata <= 8'hB4;
			14'd1201: ff_rdata <= 8'hCA;
			14'd1202: ff_rdata <= 8'hC6;
			14'd1203: ff_rdata <= 8'h44;
			14'd1204: ff_rdata <= 8'hDD;
			14'd1205: ff_rdata <= 8'h5E;
			14'd1206: ff_rdata <= 8'h04;
			14'd1207: ff_rdata <= 8'hDD;
			14'd1208: ff_rdata <= 8'h56;
			14'd1209: ff_rdata <= 8'h05;
			14'd1210: ff_rdata <= 8'h1B;
			14'd1211: ff_rdata <= 8'h7B;
			14'd1212: ff_rdata <= 8'hB2;
			14'd1213: ff_rdata <= 8'hCC;
			14'd1214: ff_rdata <= 8'hEA;
			14'd1215: ff_rdata <= 8'h44;
			14'd1216: ff_rdata <= 8'hDD;
			14'd1217: ff_rdata <= 8'h73;
			14'd1218: ff_rdata <= 8'h04;
			14'd1219: ff_rdata <= 8'hDD;
			14'd1220: ff_rdata <= 8'h72;
			14'd1221: ff_rdata <= 8'h05;
			14'd1222: ff_rdata <= 8'h11;
			14'd1223: ff_rdata <= 8'h0B;
			14'd1224: ff_rdata <= 8'h00;
			14'd1225: ff_rdata <= 8'hDD;
			14'd1226: ff_rdata <= 8'h19;
			14'd1227: ff_rdata <= 8'h10;
			14'd1228: ff_rdata <= 8'hC5;
			14'd1229: ff_rdata <= 8'hFD;
			14'd1230: ff_rdata <= 8'hE1;
			14'd1231: ff_rdata <= 8'hDD;
			14'd1232: ff_rdata <= 8'hE1;
			14'd1233: ff_rdata <= 8'hE1;
			14'd1234: ff_rdata <= 8'hD1;
			14'd1235: ff_rdata <= 8'hC1;
			14'd1236: ff_rdata <= 8'hF1;
			14'd1237: ff_rdata <= 8'hC9;
			14'd1238: ff_rdata <= 8'hDD;
			14'd1239: ff_rdata <= 8'h7E;
			14'd1240: ff_rdata <= 8'h09;
			14'd1241: ff_rdata <= 8'hB7;
			14'd1242: ff_rdata <= 8'hC0;
			14'd1243: ff_rdata <= 8'h3E;
			14'd1244: ff_rdata <= 8'h1F;
			14'd1245: ff_rdata <= 8'h80;
			14'd1246: ff_rdata <= 8'hCD;
			14'd1247: ff_rdata <= 8'h6C;
			14'd1248: ff_rdata <= 8'h41;
			14'd1249: ff_rdata <= 8'hE6;
			14'd1250: ff_rdata <= 8'hEF;
			14'd1251: ff_rdata <= 8'h5F;
			14'd1252: ff_rdata <= 8'h3E;
			14'd1253: ff_rdata <= 8'h1F;
			14'd1254: ff_rdata <= 8'h80;
			14'd1255: ff_rdata <= 8'hC3;
			14'd1256: ff_rdata <= 8'h50;
			14'd1257: ff_rdata <= 8'h41;
			14'd1258: ff_rdata <= 8'h7E;
			14'd1259: ff_rdata <= 8'h23;
			14'd1260: ff_rdata <= 8'hFE;
			14'd1261: ff_rdata <= 8'hFF;
			14'd1262: ff_rdata <= 8'hCA;
			14'd1263: ff_rdata <= 8'h24;
			14'd1264: ff_rdata <= 8'h45;
			14'd1265: ff_rdata <= 8'hFE;
			14'd1266: ff_rdata <= 8'h60;
			14'd1267: ff_rdata <= 8'hDA;
			14'd1268: ff_rdata <= 8'h54;
			14'd1269: ff_rdata <= 8'h45;
			14'd1270: ff_rdata <= 8'hFE;
			14'd1271: ff_rdata <= 8'h70;
			14'd1272: ff_rdata <= 8'hDA;
			14'd1273: ff_rdata <= 8'hDD;
			14'd1274: ff_rdata <= 8'h45;
			14'd1275: ff_rdata <= 8'hFE;
			14'd1276: ff_rdata <= 8'h80;
			14'd1277: ff_rdata <= 8'hDA;
			14'd1278: ff_rdata <= 8'hF3;
			14'd1279: ff_rdata <= 8'h45;
			14'd1280: ff_rdata <= 8'hCA;
			14'd1281: ff_rdata <= 8'h0D;
			14'd1282: ff_rdata <= 8'h46;
			14'd1283: ff_rdata <= 8'hFE;
			14'd1284: ff_rdata <= 8'h81;
			14'd1285: ff_rdata <= 8'hCA;
			14'd1286: ff_rdata <= 8'h1F;
			14'd1287: ff_rdata <= 8'h46;
			14'd1288: ff_rdata <= 8'hFE;
			14'd1289: ff_rdata <= 8'h82;
			14'd1290: ff_rdata <= 8'hCA;
			14'd1291: ff_rdata <= 8'h31;
			14'd1292: ff_rdata <= 8'h46;
			14'd1293: ff_rdata <= 8'hFE;
			14'd1294: ff_rdata <= 8'h83;
			14'd1295: ff_rdata <= 8'hCA;
			14'd1296: ff_rdata <= 8'h54;
			14'd1297: ff_rdata <= 8'h46;
			14'd1298: ff_rdata <= 8'hFE;
			14'd1299: ff_rdata <= 8'h84;
			14'd1300: ff_rdata <= 8'hCA;
			14'd1301: ff_rdata <= 8'h7A;
			14'd1302: ff_rdata <= 8'h46;
			14'd1303: ff_rdata <= 8'hFE;
			14'd1304: ff_rdata <= 8'h85;
			14'd1305: ff_rdata <= 8'hCA;
			14'd1306: ff_rdata <= 8'h73;
			14'd1307: ff_rdata <= 8'h46;
			14'd1308: ff_rdata <= 8'hFE;
			14'd1309: ff_rdata <= 8'h86;
			14'd1310: ff_rdata <= 8'hCA;
			14'd1311: ff_rdata <= 8'h6B;
			14'd1312: ff_rdata <= 8'h46;
			14'd1313: ff_rdata <= 8'hC3;
			14'd1314: ff_rdata <= 8'hEA;
			14'd1315: ff_rdata <= 8'h44;
			14'd1316: ff_rdata <= 8'hDD;
			14'd1317: ff_rdata <= 8'h36;
			14'd1318: ff_rdata <= 8'h02;
			14'd1319: ff_rdata <= 8'h00;
			14'd1320: ff_rdata <= 8'hDD;
			14'd1321: ff_rdata <= 8'h36;
			14'd1322: ff_rdata <= 8'h03;
			14'd1323: ff_rdata <= 8'h00;
			14'd1324: ff_rdata <= 8'hDD;
			14'd1325: ff_rdata <= 8'h7E;
			14'd1326: ff_rdata <= 8'h0A;
			14'd1327: ff_rdata <= 8'hB7;
			14'd1328: ff_rdata <= 8'hC8;
			14'd1329: ff_rdata <= 8'hFD;
			14'd1330: ff_rdata <= 8'h35;
			14'd1331: ff_rdata <= 8'h3C;
			14'd1332: ff_rdata <= 8'hC0;
			14'd1333: ff_rdata <= 8'hFD;
			14'd1334: ff_rdata <= 8'h7E;
			14'd1335: ff_rdata <= 8'h3A;
			14'd1336: ff_rdata <= 8'hFE;
			14'd1337: ff_rdata <= 8'hFF;
			14'd1338: ff_rdata <= 8'hCA;
			14'd1339: ff_rdata <= 8'h44;
			14'd1340: ff_rdata <= 8'h45;
			14'd1341: ff_rdata <= 8'hB7;
			14'd1342: ff_rdata <= 8'hC8;
			14'd1343: ff_rdata <= 8'h3D;
			14'd1344: ff_rdata <= 8'hFD;
			14'd1345: ff_rdata <= 8'h77;
			14'd1346: ff_rdata <= 8'h3A;
			14'd1347: ff_rdata <= 8'hC8;
			14'd1348: ff_rdata <= 8'hE1;
			14'd1349: ff_rdata <= 8'hCD;
			14'd1350: ff_rdata <= 8'h44;
			14'd1351: ff_rdata <= 8'h43;
			14'd1352: ff_rdata <= 8'hFD;
			14'd1353: ff_rdata <= 8'hE5;
			14'd1354: ff_rdata <= 8'hDD;
			14'd1355: ff_rdata <= 8'hE1;
			14'd1356: ff_rdata <= 8'h11;
			14'd1357: ff_rdata <= 8'h3D;
			14'd1358: ff_rdata <= 8'h00;
			14'd1359: ff_rdata <= 8'hDD;
			14'd1360: ff_rdata <= 8'h19;
			14'd1361: ff_rdata <= 8'hC3;
			14'd1362: ff_rdata <= 8'h65;
			14'd1363: ff_rdata <= 8'h44;
			14'd1364: ff_rdata <= 8'h4F;
			14'd1365: ff_rdata <= 8'hCD;
			14'd1366: ff_rdata <= 8'h12;
			14'd1367: ff_rdata <= 8'h47;
			14'd1368: ff_rdata <= 8'hDD;
			14'd1369: ff_rdata <= 8'h75;
			14'd1370: ff_rdata <= 8'h02;
			14'd1371: ff_rdata <= 8'hDD;
			14'd1372: ff_rdata <= 8'h74;
			14'd1373: ff_rdata <= 8'h03;
			14'd1374: ff_rdata <= 8'h79;
			14'd1375: ff_rdata <= 8'hB7;
			14'd1376: ff_rdata <= 8'hC8;
			14'd1377: ff_rdata <= 8'hD5;
			14'd1378: ff_rdata <= 8'hDD;
			14'd1379: ff_rdata <= 8'h7E;
			14'd1380: ff_rdata <= 8'h08;
			14'd1381: ff_rdata <= 8'hE6;
			14'd1382: ff_rdata <= 8'h07;
			14'd1383: ff_rdata <= 8'hC2;
			14'd1384: ff_rdata <= 8'h6F;
			14'd1385: ff_rdata <= 8'h45;
			14'd1386: ff_rdata <= 8'h63;
			14'd1387: ff_rdata <= 8'h6A;
			14'd1388: ff_rdata <= 8'hC3;
			14'd1389: ff_rdata <= 8'h8C;
			14'd1390: ff_rdata <= 8'h45;
			14'd1391: ff_rdata <= 8'h0F;
			14'd1392: ff_rdata <= 8'h0F;
			14'd1393: ff_rdata <= 8'h0F;
			14'd1394: ff_rdata <= 8'hC5;
			14'd1395: ff_rdata <= 8'h21;
			14'd1396: ff_rdata <= 8'h00;
			14'd1397: ff_rdata <= 8'h00;
			14'd1398: ff_rdata <= 8'h06;
			14'd1399: ff_rdata <= 8'h08;
			14'd1400: ff_rdata <= 8'h29;
			14'd1401: ff_rdata <= 8'h17;
			14'd1402: ff_rdata <= 8'hD2;
			14'd1403: ff_rdata <= 8'h80;
			14'd1404: ff_rdata <= 8'h45;
			14'd1405: ff_rdata <= 8'h19;
			14'd1406: ff_rdata <= 8'hCE;
			14'd1407: ff_rdata <= 8'h00;
			14'd1408: ff_rdata <= 8'h10;
			14'd1409: ff_rdata <= 8'hF6;
			14'd1410: ff_rdata <= 8'hC1;
			14'd1411: ff_rdata <= 8'h6F;
			14'd1412: ff_rdata <= 8'hB4;
			14'd1413: ff_rdata <= 8'hC2;
			14'd1414: ff_rdata <= 8'h8C;
			14'd1415: ff_rdata <= 8'h45;
			14'd1416: ff_rdata <= 8'h26;
			14'd1417: ff_rdata <= 8'h01;
			14'd1418: ff_rdata <= 8'h2E;
			14'd1419: ff_rdata <= 8'h00;
			14'd1420: ff_rdata <= 8'hDD;
			14'd1421: ff_rdata <= 8'h74;
			14'd1422: ff_rdata <= 8'h06;
			14'd1423: ff_rdata <= 8'hDD;
			14'd1424: ff_rdata <= 8'h75;
			14'd1425: ff_rdata <= 8'h07;
			14'd1426: ff_rdata <= 8'h0D;
			14'd1427: ff_rdata <= 8'h69;
			14'd1428: ff_rdata <= 8'h26;
			14'd1429: ff_rdata <= 8'h00;
			14'd1430: ff_rdata <= 8'h3E;
			14'd1431: ff_rdata <= 8'h0C;
			14'd1432: ff_rdata <= 8'hCD;
			14'd1433: ff_rdata <= 8'hC4;
			14'd1434: ff_rdata <= 8'h45;
			14'd1435: ff_rdata <= 8'h4D;
			14'd1436: ff_rdata <= 8'hCB;
			14'd1437: ff_rdata <= 8'h21;
			14'd1438: ff_rdata <= 8'h7C;
			14'd1439: ff_rdata <= 8'h87;
			14'd1440: ff_rdata <= 8'h5F;
			14'd1441: ff_rdata <= 8'h16;
			14'd1442: ff_rdata <= 8'h00;
			14'd1443: ff_rdata <= 8'h21;
			14'd1444: ff_rdata <= 8'h28;
			14'd1445: ff_rdata <= 8'h41;
			14'd1446: ff_rdata <= 8'h19;
			14'd1447: ff_rdata <= 8'h3E;
			14'd1448: ff_rdata <= 8'h0F;
			14'd1449: ff_rdata <= 8'h80;
			14'd1450: ff_rdata <= 8'h5E;
			14'd1451: ff_rdata <= 8'h23;
			14'd1452: ff_rdata <= 8'hCD;
			14'd1453: ff_rdata <= 8'h50;
			14'd1454: ff_rdata <= 8'h41;
			14'd1455: ff_rdata <= 8'h3E;
			14'd1456: ff_rdata <= 8'h1F;
			14'd1457: ff_rdata <= 8'h80;
			14'd1458: ff_rdata <= 8'hCD;
			14'd1459: ff_rdata <= 8'h6C;
			14'd1460: ff_rdata <= 8'h41;
			14'd1461: ff_rdata <= 8'hE6;
			14'd1462: ff_rdata <= 8'h20;
			14'd1463: ff_rdata <= 8'hB6;
			14'd1464: ff_rdata <= 8'hB1;
			14'd1465: ff_rdata <= 8'hF6;
			14'd1466: ff_rdata <= 8'h10;
			14'd1467: ff_rdata <= 8'h5F;
			14'd1468: ff_rdata <= 8'h3E;
			14'd1469: ff_rdata <= 8'h1F;
			14'd1470: ff_rdata <= 8'h80;
			14'd1471: ff_rdata <= 8'hCD;
			14'd1472: ff_rdata <= 8'h50;
			14'd1473: ff_rdata <= 8'h41;
			14'd1474: ff_rdata <= 8'hD1;
			14'd1475: ff_rdata <= 8'hC9;
			14'd1476: ff_rdata <= 8'hC5;
			14'd1477: ff_rdata <= 8'h06;
			14'd1478: ff_rdata <= 8'h08;
			14'd1479: ff_rdata <= 8'hB7;
			14'd1480: ff_rdata <= 8'h4F;
			14'd1481: ff_rdata <= 8'hED;
			14'd1482: ff_rdata <= 8'h6A;
			14'd1483: ff_rdata <= 8'h7C;
			14'd1484: ff_rdata <= 8'hDA;
			14'd1485: ff_rdata <= 8'hD3;
			14'd1486: ff_rdata <= 8'h45;
			14'd1487: ff_rdata <= 8'hB9;
			14'd1488: ff_rdata <= 8'hDA;
			14'd1489: ff_rdata <= 8'hD6;
			14'd1490: ff_rdata <= 8'h45;
			14'd1491: ff_rdata <= 8'h91;
			14'd1492: ff_rdata <= 8'h67;
			14'd1493: ff_rdata <= 8'hB7;
			14'd1494: ff_rdata <= 8'h3F;
			14'd1495: ff_rdata <= 8'h10;
			14'd1496: ff_rdata <= 8'hF0;
			14'd1497: ff_rdata <= 8'hCB;
			14'd1498: ff_rdata <= 8'h15;
			14'd1499: ff_rdata <= 8'hC1;
			14'd1500: ff_rdata <= 8'hC9;
			14'd1501: ff_rdata <= 8'hE6;
			14'd1502: ff_rdata <= 8'h0F;
			14'd1503: ff_rdata <= 8'h4F;
			14'd1504: ff_rdata <= 8'h3E;
			14'd1505: ff_rdata <= 8'h2F;
			14'd1506: ff_rdata <= 8'h80;
			14'd1507: ff_rdata <= 8'hCD;
			14'd1508: ff_rdata <= 8'h6C;
			14'd1509: ff_rdata <= 8'h41;
			14'd1510: ff_rdata <= 8'hE6;
			14'd1511: ff_rdata <= 8'hF0;
			14'd1512: ff_rdata <= 8'hB1;
			14'd1513: ff_rdata <= 8'h5F;
			14'd1514: ff_rdata <= 8'h3E;
			14'd1515: ff_rdata <= 8'h2F;
			14'd1516: ff_rdata <= 8'h80;
			14'd1517: ff_rdata <= 8'hCD;
			14'd1518: ff_rdata <= 8'h50;
			14'd1519: ff_rdata <= 8'h41;
			14'd1520: ff_rdata <= 8'hC3;
			14'd1521: ff_rdata <= 8'hEA;
			14'd1522: ff_rdata <= 8'h44;
			14'd1523: ff_rdata <= 8'hE6;
			14'd1524: ff_rdata <= 8'h0F;
			14'd1525: ff_rdata <= 8'h07;
			14'd1526: ff_rdata <= 8'h07;
			14'd1527: ff_rdata <= 8'h07;
			14'd1528: ff_rdata <= 8'h07;
			14'd1529: ff_rdata <= 8'h4F;
			14'd1530: ff_rdata <= 8'h3E;
			14'd1531: ff_rdata <= 8'h2F;
			14'd1532: ff_rdata <= 8'h80;
			14'd1533: ff_rdata <= 8'hCD;
			14'd1534: ff_rdata <= 8'h6C;
			14'd1535: ff_rdata <= 8'h41;
			14'd1536: ff_rdata <= 8'hE6;
			14'd1537: ff_rdata <= 8'h0F;
			14'd1538: ff_rdata <= 8'hB1;
			14'd1539: ff_rdata <= 8'h5F;
			14'd1540: ff_rdata <= 8'h3E;
			14'd1541: ff_rdata <= 8'h2F;
			14'd1542: ff_rdata <= 8'h80;
			14'd1543: ff_rdata <= 8'hCD;
			14'd1544: ff_rdata <= 8'h50;
			14'd1545: ff_rdata <= 8'h41;
			14'd1546: ff_rdata <= 8'hC3;
			14'd1547: ff_rdata <= 8'hEA;
			14'd1548: ff_rdata <= 8'h44;
			14'd1549: ff_rdata <= 8'h3E;
			14'd1550: ff_rdata <= 8'h1F;
			14'd1551: ff_rdata <= 8'h80;
			14'd1552: ff_rdata <= 8'hCD;
			14'd1553: ff_rdata <= 8'h6C;
			14'd1554: ff_rdata <= 8'h41;
			14'd1555: ff_rdata <= 8'hF6;
			14'd1556: ff_rdata <= 8'h20;
			14'd1557: ff_rdata <= 8'h5F;
			14'd1558: ff_rdata <= 8'h3E;
			14'd1559: ff_rdata <= 8'h1F;
			14'd1560: ff_rdata <= 8'h80;
			14'd1561: ff_rdata <= 8'hCD;
			14'd1562: ff_rdata <= 8'h50;
			14'd1563: ff_rdata <= 8'h41;
			14'd1564: ff_rdata <= 8'hC3;
			14'd1565: ff_rdata <= 8'hEA;
			14'd1566: ff_rdata <= 8'h44;
			14'd1567: ff_rdata <= 8'h3E;
			14'd1568: ff_rdata <= 8'h1F;
			14'd1569: ff_rdata <= 8'h80;
			14'd1570: ff_rdata <= 8'hCD;
			14'd1571: ff_rdata <= 8'h6C;
			14'd1572: ff_rdata <= 8'h41;
			14'd1573: ff_rdata <= 8'hE6;
			14'd1574: ff_rdata <= 8'hDF;
			14'd1575: ff_rdata <= 8'h5F;
			14'd1576: ff_rdata <= 8'h3E;
			14'd1577: ff_rdata <= 8'h1F;
			14'd1578: ff_rdata <= 8'h80;
			14'd1579: ff_rdata <= 8'hCD;
			14'd1580: ff_rdata <= 8'h50;
			14'd1581: ff_rdata <= 8'h41;
			14'd1582: ff_rdata <= 8'hC3;
			14'd1583: ff_rdata <= 8'hEA;
			14'd1584: ff_rdata <= 8'h44;
			14'd1585: ff_rdata <= 8'h7E;
			14'd1586: ff_rdata <= 8'h23;
			14'd1587: ff_rdata <= 8'hE6;
			14'd1588: ff_rdata <= 8'h7F;
			14'd1589: ff_rdata <= 8'hCD;
			14'd1590: ff_rdata <= 8'h3B;
			14'd1591: ff_rdata <= 8'h46;
			14'd1592: ff_rdata <= 8'hC3;
			14'd1593: ff_rdata <= 8'hEA;
			14'd1594: ff_rdata <= 8'h44;
			14'd1595: ff_rdata <= 8'h3C;
			14'd1596: ff_rdata <= 8'hE5;
			14'd1597: ff_rdata <= 8'h6F;
			14'd1598: ff_rdata <= 8'h26;
			14'd1599: ff_rdata <= 8'h00;
			14'd1600: ff_rdata <= 8'h29;
			14'd1601: ff_rdata <= 8'h29;
			14'd1602: ff_rdata <= 8'h29;
			14'd1603: ff_rdata <= 8'h11;
			14'd1604: ff_rdata <= 8'h00;
			14'd1605: ff_rdata <= 8'h4C;
			14'd1606: ff_rdata <= 8'h19;
			14'd1607: ff_rdata <= 8'h3E;
			14'd1608: ff_rdata <= 8'h07;
			14'd1609: ff_rdata <= 8'h2B;
			14'd1610: ff_rdata <= 8'h5E;
			14'd1611: ff_rdata <= 8'hCD;
			14'd1612: ff_rdata <= 8'h50;
			14'd1613: ff_rdata <= 8'h41;
			14'd1614: ff_rdata <= 8'h3D;
			14'd1615: ff_rdata <= 8'hF2;
			14'd1616: ff_rdata <= 8'h49;
			14'd1617: ff_rdata <= 8'h46;
			14'd1618: ff_rdata <= 8'hE1;
			14'd1619: ff_rdata <= 8'hC9;
			14'd1620: ff_rdata <= 8'h5E;
			14'd1621: ff_rdata <= 8'h23;
			14'd1622: ff_rdata <= 8'h56;
			14'd1623: ff_rdata <= 8'h23;
			14'd1624: ff_rdata <= 8'hE5;
			14'd1625: ff_rdata <= 8'hEB;
			14'd1626: ff_rdata <= 8'h0E;
			14'd1627: ff_rdata <= 8'h08;
			14'd1628: ff_rdata <= 8'hAF;
			14'd1629: ff_rdata <= 8'h5E;
			14'd1630: ff_rdata <= 8'h23;
			14'd1631: ff_rdata <= 8'hCD;
			14'd1632: ff_rdata <= 8'h50;
			14'd1633: ff_rdata <= 8'h41;
			14'd1634: ff_rdata <= 8'h3C;
			14'd1635: ff_rdata <= 8'h0D;
			14'd1636: ff_rdata <= 8'hC2;
			14'd1637: ff_rdata <= 8'h5D;
			14'd1638: ff_rdata <= 8'h46;
			14'd1639: ff_rdata <= 8'hE1;
			14'd1640: ff_rdata <= 8'hC3;
			14'd1641: ff_rdata <= 8'hEA;
			14'd1642: ff_rdata <= 8'h44;
			14'd1643: ff_rdata <= 8'h7E;
			14'd1644: ff_rdata <= 8'h23;
			14'd1645: ff_rdata <= 8'hDD;
			14'd1646: ff_rdata <= 8'h77;
			14'd1647: ff_rdata <= 8'h08;
			14'd1648: ff_rdata <= 8'hC3;
			14'd1649: ff_rdata <= 8'hEA;
			14'd1650: ff_rdata <= 8'h44;
			14'd1651: ff_rdata <= 8'hDD;
			14'd1652: ff_rdata <= 8'h36;
			14'd1653: ff_rdata <= 8'h09;
			14'd1654: ff_rdata <= 8'hFF;
			14'd1655: ff_rdata <= 8'hC3;
			14'd1656: ff_rdata <= 8'hEA;
			14'd1657: ff_rdata <= 8'h44;
			14'd1658: ff_rdata <= 8'hDD;
			14'd1659: ff_rdata <= 8'h36;
			14'd1660: ff_rdata <= 8'h09;
			14'd1661: ff_rdata <= 8'h00;
			14'd1662: ff_rdata <= 8'hC3;
			14'd1663: ff_rdata <= 8'hEA;
			14'd1664: ff_rdata <= 8'h44;
			14'd1665: ff_rdata <= 8'h7E;
			14'd1666: ff_rdata <= 8'h23;
			14'd1667: ff_rdata <= 8'hFE;
			14'd1668: ff_rdata <= 8'hFF;
			14'd1669: ff_rdata <= 8'hCA;
			14'd1670: ff_rdata <= 8'h24;
			14'd1671: ff_rdata <= 8'h45;
			14'd1672: ff_rdata <= 8'hB7;
			14'd1673: ff_rdata <= 8'hF2;
			14'd1674: ff_rdata <= 8'hEC;
			14'd1675: ff_rdata <= 8'h46;
			14'd1676: ff_rdata <= 8'h57;
			14'd1677: ff_rdata <= 8'h7E;
			14'd1678: ff_rdata <= 8'h23;
			14'd1679: ff_rdata <= 8'hE6;
			14'd1680: ff_rdata <= 8'h0F;
			14'd1681: ff_rdata <= 8'h4F;
			14'd1682: ff_rdata <= 8'h17;
			14'd1683: ff_rdata <= 8'h17;
			14'd1684: ff_rdata <= 8'h17;
			14'd1685: ff_rdata <= 8'h17;
			14'd1686: ff_rdata <= 8'h47;
			14'd1687: ff_rdata <= 8'hCB;
			14'd1688: ff_rdata <= 8'h1A;
			14'd1689: ff_rdata <= 8'h30;
			14'd1690: ff_rdata <= 8'h0E;
			14'd1691: ff_rdata <= 8'h3E;
			14'd1692: ff_rdata <= 8'h37;
			14'd1693: ff_rdata <= 8'hCD;
			14'd1694: ff_rdata <= 8'h6C;
			14'd1695: ff_rdata <= 8'h41;
			14'd1696: ff_rdata <= 8'hE6;
			14'd1697: ff_rdata <= 8'h0F;
			14'd1698: ff_rdata <= 8'hB0;
			14'd1699: ff_rdata <= 8'h5F;
			14'd1700: ff_rdata <= 8'h3E;
			14'd1701: ff_rdata <= 8'h37;
			14'd1702: ff_rdata <= 8'hCD;
			14'd1703: ff_rdata <= 8'h50;
			14'd1704: ff_rdata <= 8'h41;
			14'd1705: ff_rdata <= 8'hCB;
			14'd1706: ff_rdata <= 8'h1A;
			14'd1707: ff_rdata <= 8'h30;
			14'd1708: ff_rdata <= 8'h0E;
			14'd1709: ff_rdata <= 8'h3E;
			14'd1710: ff_rdata <= 8'h38;
			14'd1711: ff_rdata <= 8'hCD;
			14'd1712: ff_rdata <= 8'h6C;
			14'd1713: ff_rdata <= 8'h41;
			14'd1714: ff_rdata <= 8'hE6;
			14'd1715: ff_rdata <= 8'hF0;
			14'd1716: ff_rdata <= 8'hB1;
			14'd1717: ff_rdata <= 8'h5F;
			14'd1718: ff_rdata <= 8'h3E;
			14'd1719: ff_rdata <= 8'h38;
			14'd1720: ff_rdata <= 8'hCD;
			14'd1721: ff_rdata <= 8'h50;
			14'd1722: ff_rdata <= 8'h41;
			14'd1723: ff_rdata <= 8'hCB;
			14'd1724: ff_rdata <= 8'h1A;
			14'd1725: ff_rdata <= 8'h30;
			14'd1726: ff_rdata <= 8'h0E;
			14'd1727: ff_rdata <= 8'h3E;
			14'd1728: ff_rdata <= 8'h38;
			14'd1729: ff_rdata <= 8'hCD;
			14'd1730: ff_rdata <= 8'h6C;
			14'd1731: ff_rdata <= 8'h41;
			14'd1732: ff_rdata <= 8'hE6;
			14'd1733: ff_rdata <= 8'h0F;
			14'd1734: ff_rdata <= 8'hB0;
			14'd1735: ff_rdata <= 8'h5F;
			14'd1736: ff_rdata <= 8'h3E;
			14'd1737: ff_rdata <= 8'h38;
			14'd1738: ff_rdata <= 8'hCD;
			14'd1739: ff_rdata <= 8'h50;
			14'd1740: ff_rdata <= 8'h41;
			14'd1741: ff_rdata <= 8'hCB;
			14'd1742: ff_rdata <= 8'h1A;
			14'd1743: ff_rdata <= 8'h30;
			14'd1744: ff_rdata <= 8'h0E;
			14'd1745: ff_rdata <= 8'h3E;
			14'd1746: ff_rdata <= 8'h37;
			14'd1747: ff_rdata <= 8'hCD;
			14'd1748: ff_rdata <= 8'h6C;
			14'd1749: ff_rdata <= 8'h41;
			14'd1750: ff_rdata <= 8'hE6;
			14'd1751: ff_rdata <= 8'hF0;
			14'd1752: ff_rdata <= 8'hB1;
			14'd1753: ff_rdata <= 8'h5F;
			14'd1754: ff_rdata <= 8'h3E;
			14'd1755: ff_rdata <= 8'h37;
			14'd1756: ff_rdata <= 8'hCD;
			14'd1757: ff_rdata <= 8'h50;
			14'd1758: ff_rdata <= 8'h41;
			14'd1759: ff_rdata <= 8'hCB;
			14'd1760: ff_rdata <= 8'h1A;
			14'd1761: ff_rdata <= 8'h30;
			14'd1762: ff_rdata <= 8'h06;
			14'd1763: ff_rdata <= 8'h3E;
			14'd1764: ff_rdata <= 8'h36;
			14'd1765: ff_rdata <= 8'h59;
			14'd1766: ff_rdata <= 8'hCD;
			14'd1767: ff_rdata <= 8'h50;
			14'd1768: ff_rdata <= 8'h41;
			14'd1769: ff_rdata <= 8'hC3;
			14'd1770: ff_rdata <= 8'h81;
			14'd1771: ff_rdata <= 8'h46;
			14'd1772: ff_rdata <= 8'h4F;
			14'd1773: ff_rdata <= 8'hEE;
			14'd1774: ff_rdata <= 8'h1F;
			14'd1775: ff_rdata <= 8'h5F;
			14'd1776: ff_rdata <= 8'h3E;
			14'd1777: ff_rdata <= 8'h0E;
			14'd1778: ff_rdata <= 8'hCD;
			14'd1779: ff_rdata <= 8'h6C;
			14'd1780: ff_rdata <= 8'h41;
			14'd1781: ff_rdata <= 8'hA3;
			14'd1782: ff_rdata <= 8'h5F;
			14'd1783: ff_rdata <= 8'h3E;
			14'd1784: ff_rdata <= 8'h0E;
			14'd1785: ff_rdata <= 8'hCD;
			14'd1786: ff_rdata <= 8'h50;
			14'd1787: ff_rdata <= 8'h41;
			14'd1788: ff_rdata <= 8'hCD;
			14'd1789: ff_rdata <= 8'h6C;
			14'd1790: ff_rdata <= 8'h41;
			14'd1791: ff_rdata <= 8'h5F;
			14'd1792: ff_rdata <= 8'h79;
			14'd1793: ff_rdata <= 8'hB3;
			14'd1794: ff_rdata <= 8'h5F;
			14'd1795: ff_rdata <= 8'h3E;
			14'd1796: ff_rdata <= 8'h0E;
			14'd1797: ff_rdata <= 8'hCD;
			14'd1798: ff_rdata <= 8'h50;
			14'd1799: ff_rdata <= 8'h41;
			14'd1800: ff_rdata <= 8'hCD;
			14'd1801: ff_rdata <= 8'h12;
			14'd1802: ff_rdata <= 8'h47;
			14'd1803: ff_rdata <= 8'hDD;
			14'd1804: ff_rdata <= 8'h75;
			14'd1805: ff_rdata <= 8'h02;
			14'd1806: ff_rdata <= 8'hDD;
			14'd1807: ff_rdata <= 8'h74;
			14'd1808: ff_rdata <= 8'h03;
			14'd1809: ff_rdata <= 8'hC9;
			14'd1810: ff_rdata <= 8'h11;
			14'd1811: ff_rdata <= 8'h00;
			14'd1812: ff_rdata <= 8'h00;
			14'd1813: ff_rdata <= 8'h7E;
			14'd1814: ff_rdata <= 8'h23;
			14'd1815: ff_rdata <= 8'hFE;
			14'd1816: ff_rdata <= 8'hFF;
			14'd1817: ff_rdata <= 8'h20;
			14'd1818: ff_rdata <= 8'h04;
			14'd1819: ff_rdata <= 8'h14;
			14'd1820: ff_rdata <= 8'h1B;
			14'd1821: ff_rdata <= 8'h18;
			14'd1822: ff_rdata <= 8'hF6;
			14'd1823: ff_rdata <= 8'h83;
			14'd1824: ff_rdata <= 8'h5F;
			14'd1825: ff_rdata <= 8'h7A;
			14'd1826: ff_rdata <= 8'hCE;
			14'd1827: ff_rdata <= 8'h00;
			14'd1828: ff_rdata <= 8'h57;
			14'd1829: ff_rdata <= 8'hC9;
			14'd1830: ff_rdata <= 8'hB7;
			14'd1831: ff_rdata <= 8'hCA;
			14'd1832: ff_rdata <= 8'hDA;
			14'd1833: ff_rdata <= 8'h43;
			14'd1834: ff_rdata <= 8'h3D;
			14'd1835: ff_rdata <= 8'h87;
			14'd1836: ff_rdata <= 8'h16;
			14'd1837: ff_rdata <= 8'h00;
			14'd1838: ff_rdata <= 8'h5F;
			14'd1839: ff_rdata <= 8'h21;
			14'd1840: ff_rdata <= 8'h10;
			14'd1841: ff_rdata <= 8'h80;
			14'd1842: ff_rdata <= 8'h19;
			14'd1843: ff_rdata <= 8'h7E;
			14'd1844: ff_rdata <= 8'h23;
			14'd1845: ff_rdata <= 8'h66;
			14'd1846: ff_rdata <= 8'h6F;
			14'd1847: ff_rdata <= 8'h78;
			14'd1848: ff_rdata <= 8'hC3;
			14'd1849: ff_rdata <= 8'hCE;
			14'd1850: ff_rdata <= 8'h42;
			14'd1851: ff_rdata <= 8'hC5;
			14'd1852: ff_rdata <= 8'hE5;
			14'd1853: ff_rdata <= 8'h01;
			14'd1854: ff_rdata <= 8'h00;
			14'd1855: ff_rdata <= 8'h40;
			14'd1856: ff_rdata <= 8'hCD;
			14'd1857: ff_rdata <= 8'hDC;
			14'd1858: ff_rdata <= 8'h41;
			14'd1859: ff_rdata <= 8'h7E;
			14'd1860: ff_rdata <= 8'h23;
			14'd1861: ff_rdata <= 8'h66;
			14'd1862: ff_rdata <= 8'hE6;
			14'd1863: ff_rdata <= 8'hFE;
			14'd1864: ff_rdata <= 8'h6F;
			14'd1865: ff_rdata <= 8'h01;
			14'd1866: ff_rdata <= 8'h3A;
			14'd1867: ff_rdata <= 8'h00;
			14'd1868: ff_rdata <= 8'h09;
			14'd1869: ff_rdata <= 8'h7E;
			14'd1870: ff_rdata <= 8'hE1;
			14'd1871: ff_rdata <= 8'hC1;
			14'd1872: ff_rdata <= 8'hC9;
			14'd1873: ff_rdata <= 8'h00;
			14'd1874: ff_rdata <= 8'h00;
			14'd1875: ff_rdata <= 8'hE1;
			14'd1876: ff_rdata <= 8'h00;
			14'd1877: ff_rdata <= 8'h00;
			14'd1878: ff_rdata <= 8'h00;
			14'd1879: ff_rdata <= 8'h00;
			14'd1880: ff_rdata <= 8'h00;
			14'd1881: ff_rdata <= 8'h00;
			14'd1882: ff_rdata <= 8'h00;
			14'd1883: ff_rdata <= 8'h00;
			14'd1884: ff_rdata <= 8'h00;
			14'd1885: ff_rdata <= 8'h00;
			14'd1886: ff_rdata <= 8'h00;
			14'd1887: ff_rdata <= 8'h00;
			14'd1888: ff_rdata <= 8'h00;
			14'd1889: ff_rdata <= 8'h00;
			14'd1890: ff_rdata <= 8'h00;
			14'd1891: ff_rdata <= 8'h00;
			14'd1892: ff_rdata <= 8'h00;
			14'd1893: ff_rdata <= 8'h00;
			14'd1894: ff_rdata <= 8'h00;
			14'd1895: ff_rdata <= 8'h00;
			14'd1896: ff_rdata <= 8'h00;
			14'd1897: ff_rdata <= 8'h00;
			14'd1898: ff_rdata <= 8'h00;
			14'd1899: ff_rdata <= 8'h00;
			14'd1900: ff_rdata <= 8'hE4;
			14'd1901: ff_rdata <= 8'h00;
			14'd1902: ff_rdata <= 8'h00;
			14'd1903: ff_rdata <= 8'h00;
			14'd1904: ff_rdata <= 8'h00;
			14'd1905: ff_rdata <= 8'h00;
			14'd1906: ff_rdata <= 8'h00;
			14'd1907: ff_rdata <= 8'h00;
			14'd1908: ff_rdata <= 8'h00;
			14'd1909: ff_rdata <= 8'h00;
			14'd1910: ff_rdata <= 8'h00;
			14'd1911: ff_rdata <= 8'h00;
			14'd1912: ff_rdata <= 8'h00;
			14'd1913: ff_rdata <= 8'h00;
			14'd1914: ff_rdata <= 8'h00;
			14'd1915: ff_rdata <= 8'h00;
			14'd1916: ff_rdata <= 8'h00;
			14'd1917: ff_rdata <= 8'h00;
			14'd1918: ff_rdata <= 8'h00;
			14'd1919: ff_rdata <= 8'h8A;
			14'd1920: ff_rdata <= 8'hDE;
			14'd1921: ff_rdata <= 8'hFF;
			14'd1922: ff_rdata <= 8'hFF;
			14'd1923: ff_rdata <= 8'hFF;
			14'd1924: ff_rdata <= 8'hFF;
			14'd1925: ff_rdata <= 8'hE7;
			14'd1926: ff_rdata <= 8'hFF;
			14'd1927: ff_rdata <= 8'hFF;
			14'd1928: ff_rdata <= 8'hFF;
			14'd1929: ff_rdata <= 8'hFF;
			14'd1930: ff_rdata <= 8'hFF;
			14'd1931: ff_rdata <= 8'hFF;
			14'd1932: ff_rdata <= 8'hFF;
			14'd1933: ff_rdata <= 8'hFF;
			14'd1934: ff_rdata <= 8'hFF;
			14'd1935: ff_rdata <= 8'hFF;
			14'd1936: ff_rdata <= 8'hFF;
			14'd1937: ff_rdata <= 8'hFF;
			14'd1938: ff_rdata <= 8'hFF;
			14'd1939: ff_rdata <= 8'hFF;
			14'd1940: ff_rdata <= 8'hFF;
			14'd1941: ff_rdata <= 8'hFF;
			14'd1942: ff_rdata <= 8'hFF;
			14'd1943: ff_rdata <= 8'hFF;
			14'd1944: ff_rdata <= 8'hFF;
			14'd1945: ff_rdata <= 8'hFF;
			14'd1946: ff_rdata <= 8'hFF;
			14'd1947: ff_rdata <= 8'hFF;
			14'd1948: ff_rdata <= 8'hFF;
			14'd1949: ff_rdata <= 8'hFF;
			14'd1950: ff_rdata <= 8'hEA;
			14'd1951: ff_rdata <= 8'hFF;
			14'd1952: ff_rdata <= 8'hFF;
			14'd1953: ff_rdata <= 8'hFF;
			14'd1954: ff_rdata <= 8'hFF;
			14'd1955: ff_rdata <= 8'hFF;
			14'd1956: ff_rdata <= 8'hFF;
			14'd1957: ff_rdata <= 8'hFF;
			14'd1958: ff_rdata <= 8'hFF;
			14'd1959: ff_rdata <= 8'hFF;
			14'd1960: ff_rdata <= 8'hFF;
			14'd1961: ff_rdata <= 8'hFF;
			14'd1962: ff_rdata <= 8'hFF;
			14'd1963: ff_rdata <= 8'hFF;
			14'd1964: ff_rdata <= 8'hFF;
			14'd1965: ff_rdata <= 8'hFF;
			14'd1966: ff_rdata <= 8'hFF;
			14'd1967: ff_rdata <= 8'hFF;
			14'd1968: ff_rdata <= 8'hFF;
			14'd1969: ff_rdata <= 8'hFF;
			14'd1970: ff_rdata <= 8'hFF;
			14'd1971: ff_rdata <= 8'hFF;
			14'd1972: ff_rdata <= 8'hFF;
			14'd1973: ff_rdata <= 8'hFF;
			14'd1974: ff_rdata <= 8'hFF;
			14'd1975: ff_rdata <= 8'hED;
			14'd1976: ff_rdata <= 8'hFF;
			14'd1977: ff_rdata <= 8'hFF;
			14'd1978: ff_rdata <= 8'hFF;
			14'd1979: ff_rdata <= 8'hFF;
			14'd1980: ff_rdata <= 8'hFF;
			14'd1981: ff_rdata <= 8'hFF;
			14'd1982: ff_rdata <= 8'hFF;
			14'd1983: ff_rdata <= 8'hFF;
			14'd1984: ff_rdata <= 8'h00;
			14'd1985: ff_rdata <= 8'h00;
			14'd1986: ff_rdata <= 8'h00;
			14'd1987: ff_rdata <= 8'h00;
			14'd1988: ff_rdata <= 8'h00;
			14'd1989: ff_rdata <= 8'h00;
			14'd1990: ff_rdata <= 8'h00;
			14'd1991: ff_rdata <= 8'h00;
			14'd1992: ff_rdata <= 8'h00;
			14'd1993: ff_rdata <= 8'h00;
			14'd1994: ff_rdata <= 8'h00;
			14'd1995: ff_rdata <= 8'h00;
			14'd1996: ff_rdata <= 8'h00;
			14'd1997: ff_rdata <= 8'h00;
			14'd1998: ff_rdata <= 8'h00;
			14'd1999: ff_rdata <= 8'h00;
			14'd2000: ff_rdata <= 8'hF0;
			14'd2001: ff_rdata <= 8'h00;
			14'd2002: ff_rdata <= 8'h00;
			14'd2003: ff_rdata <= 8'h00;
			14'd2004: ff_rdata <= 8'h00;
			14'd2005: ff_rdata <= 8'h00;
			14'd2006: ff_rdata <= 8'h00;
			14'd2007: ff_rdata <= 8'h00;
			14'd2008: ff_rdata <= 8'h00;
			14'd2009: ff_rdata <= 8'h00;
			14'd2010: ff_rdata <= 8'h00;
			14'd2011: ff_rdata <= 8'h00;
			14'd2012: ff_rdata <= 8'h00;
			14'd2013: ff_rdata <= 8'h00;
			14'd2014: ff_rdata <= 8'h00;
			14'd2015: ff_rdata <= 8'h00;
			14'd2016: ff_rdata <= 8'h00;
			14'd2017: ff_rdata <= 8'h00;
			14'd2018: ff_rdata <= 8'h00;
			14'd2019: ff_rdata <= 8'h00;
			14'd2020: ff_rdata <= 8'h00;
			14'd2021: ff_rdata <= 8'h00;
			14'd2022: ff_rdata <= 8'h00;
			14'd2023: ff_rdata <= 8'h00;
			14'd2024: ff_rdata <= 8'h00;
			14'd2025: ff_rdata <= 8'hF3;
			14'd2026: ff_rdata <= 8'h00;
			14'd2027: ff_rdata <= 8'h00;
			14'd2028: ff_rdata <= 8'h00;
			14'd2029: ff_rdata <= 8'h00;
			14'd2030: ff_rdata <= 8'h00;
			14'd2031: ff_rdata <= 8'h00;
			14'd2032: ff_rdata <= 8'h00;
			14'd2033: ff_rdata <= 8'h00;
			14'd2034: ff_rdata <= 8'h00;
			14'd2035: ff_rdata <= 8'h00;
			14'd2036: ff_rdata <= 8'h00;
			14'd2037: ff_rdata <= 8'h00;
			14'd2038: ff_rdata <= 8'h00;
			14'd2039: ff_rdata <= 8'h00;
			14'd2040: ff_rdata <= 8'h00;
			14'd2041: ff_rdata <= 8'h00;
			14'd2042: ff_rdata <= 8'h00;
			14'd2043: ff_rdata <= 8'h00;
			14'd2044: ff_rdata <= 8'h00;
			14'd2045: ff_rdata <= 8'h00;
			14'd2046: ff_rdata <= 8'h00;
			14'd2047: ff_rdata <= 8'h00;
			14'd2048: ff_rdata <= 8'hFF;
			14'd2049: ff_rdata <= 8'hFF;
			14'd2050: ff_rdata <= 8'hF6;
			14'd2051: ff_rdata <= 8'hFF;
			14'd2052: ff_rdata <= 8'hFF;
			14'd2053: ff_rdata <= 8'hFF;
			14'd2054: ff_rdata <= 8'hFF;
			14'd2055: ff_rdata <= 8'hFF;
			14'd2056: ff_rdata <= 8'hFF;
			14'd2057: ff_rdata <= 8'hFF;
			14'd2058: ff_rdata <= 8'hFF;
			14'd2059: ff_rdata <= 8'hFF;
			14'd2060: ff_rdata <= 8'hFF;
			14'd2061: ff_rdata <= 8'hFF;
			14'd2062: ff_rdata <= 8'hFF;
			14'd2063: ff_rdata <= 8'hFF;
			14'd2064: ff_rdata <= 8'hFF;
			14'd2065: ff_rdata <= 8'hFF;
			14'd2066: ff_rdata <= 8'hFF;
			14'd2067: ff_rdata <= 8'hFF;
			14'd2068: ff_rdata <= 8'hFF;
			14'd2069: ff_rdata <= 8'hFF;
			14'd2070: ff_rdata <= 8'hFF;
			14'd2071: ff_rdata <= 8'hFF;
			14'd2072: ff_rdata <= 8'hFF;
			14'd2073: ff_rdata <= 8'hFF;
			14'd2074: ff_rdata <= 8'hFF;
			14'd2075: ff_rdata <= 8'hF9;
			14'd2076: ff_rdata <= 8'hFF;
			14'd2077: ff_rdata <= 8'hFF;
			14'd2078: ff_rdata <= 8'hFF;
			14'd2079: ff_rdata <= 8'hFF;
			14'd2080: ff_rdata <= 8'hFF;
			14'd2081: ff_rdata <= 8'hFF;
			14'd2082: ff_rdata <= 8'hFF;
			14'd2083: ff_rdata <= 8'hFF;
			14'd2084: ff_rdata <= 8'hFF;
			14'd2085: ff_rdata <= 8'hFF;
			14'd2086: ff_rdata <= 8'hFF;
			14'd2087: ff_rdata <= 8'hFF;
			14'd2088: ff_rdata <= 8'hFF;
			14'd2089: ff_rdata <= 8'hFF;
			14'd2090: ff_rdata <= 8'hFF;
			14'd2091: ff_rdata <= 8'hFF;
			14'd2092: ff_rdata <= 8'hFF;
			14'd2093: ff_rdata <= 8'hFF;
			14'd2094: ff_rdata <= 8'hFF;
			14'd2095: ff_rdata <= 8'hFF;
			14'd2096: ff_rdata <= 8'hFF;
			14'd2097: ff_rdata <= 8'hFF;
			14'd2098: ff_rdata <= 8'hFF;
			14'd2099: ff_rdata <= 8'hFF;
			14'd2100: ff_rdata <= 8'hFC;
			14'd2101: ff_rdata <= 8'hFF;
			14'd2102: ff_rdata <= 8'hFF;
			14'd2103: ff_rdata <= 8'hFF;
			14'd2104: ff_rdata <= 8'hFF;
			14'd2105: ff_rdata <= 8'hFF;
			14'd2106: ff_rdata <= 8'hFF;
			14'd2107: ff_rdata <= 8'hFF;
			14'd2108: ff_rdata <= 8'hFF;
			14'd2109: ff_rdata <= 8'hFF;
			14'd2110: ff_rdata <= 8'hFF;
			14'd2111: ff_rdata <= 8'hFF;
			14'd2112: ff_rdata <= 8'h00;
			14'd2113: ff_rdata <= 8'h00;
			14'd2114: ff_rdata <= 8'h00;
			14'd2115: ff_rdata <= 8'h00;
			14'd2116: ff_rdata <= 8'h00;
			14'd2117: ff_rdata <= 8'h00;
			14'd2118: ff_rdata <= 8'h00;
			14'd2119: ff_rdata <= 8'h00;
			14'd2120: ff_rdata <= 8'h00;
			14'd2121: ff_rdata <= 8'h00;
			14'd2122: ff_rdata <= 8'h00;
			14'd2123: ff_rdata <= 8'h00;
			14'd2124: ff_rdata <= 8'h00;
			14'd2125: ff_rdata <= 8'hFF;
			14'd2126: ff_rdata <= 8'h00;
			14'd2127: ff_rdata <= 8'h00;
			14'd2128: ff_rdata <= 8'h00;
			14'd2129: ff_rdata <= 8'h00;
			14'd2130: ff_rdata <= 8'h00;
			14'd2131: ff_rdata <= 8'h00;
			14'd2132: ff_rdata <= 8'h00;
			14'd2133: ff_rdata <= 8'h00;
			14'd2134: ff_rdata <= 8'h00;
			14'd2135: ff_rdata <= 8'h00;
			14'd2136: ff_rdata <= 8'h00;
			14'd2137: ff_rdata <= 8'h00;
			14'd2138: ff_rdata <= 8'h00;
			14'd2139: ff_rdata <= 8'h00;
			14'd2140: ff_rdata <= 8'h00;
			14'd2141: ff_rdata <= 8'h00;
			14'd2142: ff_rdata <= 8'h00;
			14'd2143: ff_rdata <= 8'h00;
			14'd2144: ff_rdata <= 8'h00;
			14'd2145: ff_rdata <= 8'h00;
			14'd2146: ff_rdata <= 8'h00;
			14'd2147: ff_rdata <= 8'h00;
			14'd2148: ff_rdata <= 8'h00;
			14'd2149: ff_rdata <= 8'h00;
			14'd2150: ff_rdata <= 8'h02;
			14'd2151: ff_rdata <= 8'h00;
			14'd2152: ff_rdata <= 8'h00;
			14'd2153: ff_rdata <= 8'h00;
			14'd2154: ff_rdata <= 8'h00;
			14'd2155: ff_rdata <= 8'h00;
			14'd2156: ff_rdata <= 8'h00;
			14'd2157: ff_rdata <= 8'h00;
			14'd2158: ff_rdata <= 8'h00;
			14'd2159: ff_rdata <= 8'h00;
			14'd2160: ff_rdata <= 8'h00;
			14'd2161: ff_rdata <= 8'h00;
			14'd2162: ff_rdata <= 8'h00;
			14'd2163: ff_rdata <= 8'h00;
			14'd2164: ff_rdata <= 8'h00;
			14'd2165: ff_rdata <= 8'h00;
			14'd2166: ff_rdata <= 8'h00;
			14'd2167: ff_rdata <= 8'h00;
			14'd2168: ff_rdata <= 8'h00;
			14'd2169: ff_rdata <= 8'h00;
			14'd2170: ff_rdata <= 8'h00;
			14'd2171: ff_rdata <= 8'h00;
			14'd2172: ff_rdata <= 8'h00;
			14'd2173: ff_rdata <= 8'h00;
			14'd2174: ff_rdata <= 8'h00;
			14'd2175: ff_rdata <= 8'h05;
			14'd2176: ff_rdata <= 8'hDF;
			14'd2177: ff_rdata <= 8'hFF;
			14'd2178: ff_rdata <= 8'hFF;
			14'd2179: ff_rdata <= 8'hFF;
			14'd2180: ff_rdata <= 8'hFF;
			14'd2181: ff_rdata <= 8'hFF;
			14'd2182: ff_rdata <= 8'hFF;
			14'd2183: ff_rdata <= 8'hFF;
			14'd2184: ff_rdata <= 8'hFF;
			14'd2185: ff_rdata <= 8'hFF;
			14'd2186: ff_rdata <= 8'hFF;
			14'd2187: ff_rdata <= 8'hFF;
			14'd2188: ff_rdata <= 8'hFF;
			14'd2189: ff_rdata <= 8'hFF;
			14'd2190: ff_rdata <= 8'hFF;
			14'd2191: ff_rdata <= 8'hFF;
			14'd2192: ff_rdata <= 8'hFF;
			14'd2193: ff_rdata <= 8'hFF;
			14'd2194: ff_rdata <= 8'hFF;
			14'd2195: ff_rdata <= 8'hFF;
			14'd2196: ff_rdata <= 8'hFF;
			14'd2197: ff_rdata <= 8'hFF;
			14'd2198: ff_rdata <= 8'hFF;
			14'd2199: ff_rdata <= 8'hFF;
			14'd2200: ff_rdata <= 8'h08;
			14'd2201: ff_rdata <= 8'hFF;
			14'd2202: ff_rdata <= 8'hFF;
			14'd2203: ff_rdata <= 8'hFF;
			14'd2204: ff_rdata <= 8'hFF;
			14'd2205: ff_rdata <= 8'hFF;
			14'd2206: ff_rdata <= 8'hFF;
			14'd2207: ff_rdata <= 8'hFF;
			14'd2208: ff_rdata <= 8'hFF;
			14'd2209: ff_rdata <= 8'hFF;
			14'd2210: ff_rdata <= 8'hFF;
			14'd2211: ff_rdata <= 8'hFF;
			14'd2212: ff_rdata <= 8'hFF;
			14'd2213: ff_rdata <= 8'hFF;
			14'd2214: ff_rdata <= 8'hFF;
			14'd2215: ff_rdata <= 8'hFF;
			14'd2216: ff_rdata <= 8'hFF;
			14'd2217: ff_rdata <= 8'hFF;
			14'd2218: ff_rdata <= 8'hFF;
			14'd2219: ff_rdata <= 8'hFF;
			14'd2220: ff_rdata <= 8'hFF;
			14'd2221: ff_rdata <= 8'hFF;
			14'd2222: ff_rdata <= 8'hFF;
			14'd2223: ff_rdata <= 8'hFF;
			14'd2224: ff_rdata <= 8'hFF;
			14'd2225: ff_rdata <= 8'h0B;
			14'd2226: ff_rdata <= 8'hFF;
			14'd2227: ff_rdata <= 8'hFF;
			14'd2228: ff_rdata <= 8'hFF;
			14'd2229: ff_rdata <= 8'hFF;
			14'd2230: ff_rdata <= 8'hFF;
			14'd2231: ff_rdata <= 8'hFF;
			14'd2232: ff_rdata <= 8'hFF;
			14'd2233: ff_rdata <= 8'hFF;
			14'd2234: ff_rdata <= 8'hFF;
			14'd2235: ff_rdata <= 8'hFF;
			14'd2236: ff_rdata <= 8'hFF;
			14'd2237: ff_rdata <= 8'hFF;
			14'd2238: ff_rdata <= 8'hFF;
			14'd2239: ff_rdata <= 8'hFF;
			14'd2240: ff_rdata <= 8'h00;
			14'd2241: ff_rdata <= 8'h00;
			14'd2242: ff_rdata <= 8'h00;
			14'd2243: ff_rdata <= 8'h00;
			14'd2244: ff_rdata <= 8'h00;
			14'd2245: ff_rdata <= 8'h00;
			14'd2246: ff_rdata <= 8'h00;
			14'd2247: ff_rdata <= 8'h00;
			14'd2248: ff_rdata <= 8'h00;
			14'd2249: ff_rdata <= 8'h00;
			14'd2250: ff_rdata <= 8'h0E;
			14'd2251: ff_rdata <= 8'h00;
			14'd2252: ff_rdata <= 8'h00;
			14'd2253: ff_rdata <= 8'h00;
			14'd2254: ff_rdata <= 8'h00;
			14'd2255: ff_rdata <= 8'h00;
			14'd2256: ff_rdata <= 8'h00;
			14'd2257: ff_rdata <= 8'h00;
			14'd2258: ff_rdata <= 8'h00;
			14'd2259: ff_rdata <= 8'h00;
			14'd2260: ff_rdata <= 8'h00;
			14'd2261: ff_rdata <= 8'h00;
			14'd2262: ff_rdata <= 8'h00;
			14'd2263: ff_rdata <= 8'h00;
			14'd2264: ff_rdata <= 8'h00;
			14'd2265: ff_rdata <= 8'h00;
			14'd2266: ff_rdata <= 8'h00;
			14'd2267: ff_rdata <= 8'h00;
			14'd2268: ff_rdata <= 8'h00;
			14'd2269: ff_rdata <= 8'h00;
			14'd2270: ff_rdata <= 8'h00;
			14'd2271: ff_rdata <= 8'h00;
			14'd2272: ff_rdata <= 8'h00;
			14'd2273: ff_rdata <= 8'h00;
			14'd2274: ff_rdata <= 8'h00;
			14'd2275: ff_rdata <= 8'h11;
			14'd2276: ff_rdata <= 8'h00;
			14'd2277: ff_rdata <= 8'h00;
			14'd2278: ff_rdata <= 8'h00;
			14'd2279: ff_rdata <= 8'h00;
			14'd2280: ff_rdata <= 8'h00;
			14'd2281: ff_rdata <= 8'h00;
			14'd2282: ff_rdata <= 8'h00;
			14'd2283: ff_rdata <= 8'h00;
			14'd2284: ff_rdata <= 8'h00;
			14'd2285: ff_rdata <= 8'h00;
			14'd2286: ff_rdata <= 8'h00;
			14'd2287: ff_rdata <= 8'h00;
			14'd2288: ff_rdata <= 8'h00;
			14'd2289: ff_rdata <= 8'h00;
			14'd2290: ff_rdata <= 8'h00;
			14'd2291: ff_rdata <= 8'h00;
			14'd2292: ff_rdata <= 8'h00;
			14'd2293: ff_rdata <= 8'h00;
			14'd2294: ff_rdata <= 8'h00;
			14'd2295: ff_rdata <= 8'h00;
			14'd2296: ff_rdata <= 8'h00;
			14'd2297: ff_rdata <= 8'h00;
			14'd2298: ff_rdata <= 8'h00;
			14'd2299: ff_rdata <= 8'h00;
			14'd2300: ff_rdata <= 8'h14;
			14'd2301: ff_rdata <= 8'h00;
			14'd2302: ff_rdata <= 8'h00;
			14'd2303: ff_rdata <= 8'h0E;
			14'd2304: ff_rdata <= 8'h00;
			14'd2305: ff_rdata <= 8'h00;
			14'd2306: ff_rdata <= 8'h00;
			14'd2307: ff_rdata <= 8'h00;
			14'd2308: ff_rdata <= 8'h00;
			14'd2309: ff_rdata <= 8'h00;
			14'd2310: ff_rdata <= 8'h00;
			14'd2311: ff_rdata <= 8'h00;
			14'd2312: ff_rdata <= 8'h00;
			14'd2313: ff_rdata <= 8'h00;
			14'd2314: ff_rdata <= 8'h00;
			14'd2315: ff_rdata <= 8'h00;
			14'd2316: ff_rdata <= 8'h00;
			14'd2317: ff_rdata <= 8'h00;
			14'd2318: ff_rdata <= 8'h00;
			14'd2319: ff_rdata <= 8'h00;
			14'd2320: ff_rdata <= 8'h00;
			14'd2321: ff_rdata <= 8'h00;
			14'd2322: ff_rdata <= 8'h00;
			14'd2323: ff_rdata <= 8'h00;
			14'd2324: ff_rdata <= 8'h00;
			14'd2325: ff_rdata <= 8'h17;
			14'd2326: ff_rdata <= 8'h00;
			14'd2327: ff_rdata <= 8'h00;
			14'd2328: ff_rdata <= 8'h00;
			14'd2329: ff_rdata <= 8'h00;
			14'd2330: ff_rdata <= 8'h00;
			14'd2331: ff_rdata <= 8'h00;
			14'd2332: ff_rdata <= 8'h00;
			14'd2333: ff_rdata <= 8'h00;
			14'd2334: ff_rdata <= 8'h00;
			14'd2335: ff_rdata <= 8'h00;
			14'd2336: ff_rdata <= 8'h00;
			14'd2337: ff_rdata <= 8'h00;
			14'd2338: ff_rdata <= 8'h00;
			14'd2339: ff_rdata <= 8'h00;
			14'd2340: ff_rdata <= 8'h00;
			14'd2341: ff_rdata <= 8'h00;
			14'd2342: ff_rdata <= 8'h00;
			14'd2343: ff_rdata <= 8'h00;
			14'd2344: ff_rdata <= 8'h00;
			14'd2345: ff_rdata <= 8'h00;
			14'd2346: ff_rdata <= 8'h00;
			14'd2347: ff_rdata <= 8'h00;
			14'd2348: ff_rdata <= 8'h00;
			14'd2349: ff_rdata <= 8'h00;
			14'd2350: ff_rdata <= 8'h1A;
			14'd2351: ff_rdata <= 8'h00;
			14'd2352: ff_rdata <= 8'h00;
			14'd2353: ff_rdata <= 8'h00;
			14'd2354: ff_rdata <= 8'h00;
			14'd2355: ff_rdata <= 8'h00;
			14'd2356: ff_rdata <= 8'h00;
			14'd2357: ff_rdata <= 8'h00;
			14'd2358: ff_rdata <= 8'h00;
			14'd2359: ff_rdata <= 8'h00;
			14'd2360: ff_rdata <= 8'h00;
			14'd2361: ff_rdata <= 8'h00;
			14'd2362: ff_rdata <= 8'h00;
			14'd2363: ff_rdata <= 8'h00;
			14'd2364: ff_rdata <= 8'h00;
			14'd2365: ff_rdata <= 8'h00;
			14'd2366: ff_rdata <= 8'h00;
			14'd2367: ff_rdata <= 8'h00;
			14'd2368: ff_rdata <= 8'hFF;
			14'd2369: ff_rdata <= 8'hFF;
			14'd2370: ff_rdata <= 8'hFF;
			14'd2371: ff_rdata <= 8'hFF;
			14'd2372: ff_rdata <= 8'hFF;
			14'd2373: ff_rdata <= 8'hFF;
			14'd2374: ff_rdata <= 8'hFF;
			14'd2375: ff_rdata <= 8'h1D;
			14'd2376: ff_rdata <= 8'hFF;
			14'd2377: ff_rdata <= 8'hFF;
			14'd2378: ff_rdata <= 8'hFF;
			14'd2379: ff_rdata <= 8'hFF;
			14'd2380: ff_rdata <= 8'hFF;
			14'd2381: ff_rdata <= 8'hFF;
			14'd2382: ff_rdata <= 8'hFF;
			14'd2383: ff_rdata <= 8'hFF;
			14'd2384: ff_rdata <= 8'hFF;
			14'd2385: ff_rdata <= 8'hFF;
			14'd2386: ff_rdata <= 8'hFF;
			14'd2387: ff_rdata <= 8'hFF;
			14'd2388: ff_rdata <= 8'hFF;
			14'd2389: ff_rdata <= 8'hFF;
			14'd2390: ff_rdata <= 8'hFF;
			14'd2391: ff_rdata <= 8'hFF;
			14'd2392: ff_rdata <= 8'hFF;
			14'd2393: ff_rdata <= 8'hFF;
			14'd2394: ff_rdata <= 8'hFF;
			14'd2395: ff_rdata <= 8'hFF;
			14'd2396: ff_rdata <= 8'hFF;
			14'd2397: ff_rdata <= 8'hFF;
			14'd2398: ff_rdata <= 8'hFF;
			14'd2399: ff_rdata <= 8'hFF;
			14'd2400: ff_rdata <= 8'h20;
			14'd2401: ff_rdata <= 8'hFF;
			14'd2402: ff_rdata <= 8'hFF;
			14'd2403: ff_rdata <= 8'hFF;
			14'd2404: ff_rdata <= 8'hFF;
			14'd2405: ff_rdata <= 8'hFF;
			14'd2406: ff_rdata <= 8'hFF;
			14'd2407: ff_rdata <= 8'hFF;
			14'd2408: ff_rdata <= 8'hFF;
			14'd2409: ff_rdata <= 8'hFF;
			14'd2410: ff_rdata <= 8'hFF;
			14'd2411: ff_rdata <= 8'hFF;
			14'd2412: ff_rdata <= 8'hFF;
			14'd2413: ff_rdata <= 8'hFF;
			14'd2414: ff_rdata <= 8'hFF;
			14'd2415: ff_rdata <= 8'hFF;
			14'd2416: ff_rdata <= 8'hFF;
			14'd2417: ff_rdata <= 8'hFF;
			14'd2418: ff_rdata <= 8'hFF;
			14'd2419: ff_rdata <= 8'hFF;
			14'd2420: ff_rdata <= 8'hFF;
			14'd2421: ff_rdata <= 8'hFF;
			14'd2422: ff_rdata <= 8'hFF;
			14'd2423: ff_rdata <= 8'hFF;
			14'd2424: ff_rdata <= 8'hFF;
			14'd2425: ff_rdata <= 8'h23;
			14'd2426: ff_rdata <= 8'hFF;
			14'd2427: ff_rdata <= 8'hFF;
			14'd2428: ff_rdata <= 8'hFF;
			14'd2429: ff_rdata <= 8'hFF;
			14'd2430: ff_rdata <= 8'hFF;
			14'd2431: ff_rdata <= 8'h37;
			14'd2432: ff_rdata <= 8'h21;
			14'd2433: ff_rdata <= 8'h00;
			14'd2434: ff_rdata <= 8'h00;
			14'd2435: ff_rdata <= 8'h00;
			14'd2436: ff_rdata <= 8'h00;
			14'd2437: ff_rdata <= 8'h00;
			14'd2438: ff_rdata <= 8'h00;
			14'd2439: ff_rdata <= 8'h00;
			14'd2440: ff_rdata <= 8'h00;
			14'd2441: ff_rdata <= 8'h00;
			14'd2442: ff_rdata <= 8'h00;
			14'd2443: ff_rdata <= 8'h00;
			14'd2444: ff_rdata <= 8'h00;
			14'd2445: ff_rdata <= 8'h00;
			14'd2446: ff_rdata <= 8'h00;
			14'd2447: ff_rdata <= 8'h00;
			14'd2448: ff_rdata <= 8'h00;
			14'd2449: ff_rdata <= 8'h00;
			14'd2450: ff_rdata <= 8'h26;
			14'd2451: ff_rdata <= 8'h00;
			14'd2452: ff_rdata <= 8'h00;
			14'd2453: ff_rdata <= 8'h00;
			14'd2454: ff_rdata <= 8'h00;
			14'd2455: ff_rdata <= 8'h00;
			14'd2456: ff_rdata <= 8'h00;
			14'd2457: ff_rdata <= 8'h00;
			14'd2458: ff_rdata <= 8'h00;
			14'd2459: ff_rdata <= 8'h00;
			14'd2460: ff_rdata <= 8'h00;
			14'd2461: ff_rdata <= 8'h00;
			14'd2462: ff_rdata <= 8'h00;
			14'd2463: ff_rdata <= 8'h00;
			14'd2464: ff_rdata <= 8'h00;
			14'd2465: ff_rdata <= 8'h00;
			14'd2466: ff_rdata <= 8'h00;
			14'd2467: ff_rdata <= 8'h00;
			14'd2468: ff_rdata <= 8'h00;
			14'd2469: ff_rdata <= 8'h00;
			14'd2470: ff_rdata <= 8'h00;
			14'd2471: ff_rdata <= 8'h00;
			14'd2472: ff_rdata <= 8'h00;
			14'd2473: ff_rdata <= 8'h00;
			14'd2474: ff_rdata <= 8'h00;
			14'd2475: ff_rdata <= 8'h29;
			14'd2476: ff_rdata <= 8'h00;
			14'd2477: ff_rdata <= 8'h00;
			14'd2478: ff_rdata <= 8'h00;
			14'd2479: ff_rdata <= 8'h00;
			14'd2480: ff_rdata <= 8'h00;
			14'd2481: ff_rdata <= 8'h00;
			14'd2482: ff_rdata <= 8'h00;
			14'd2483: ff_rdata <= 8'h00;
			14'd2484: ff_rdata <= 8'h00;
			14'd2485: ff_rdata <= 8'h00;
			14'd2486: ff_rdata <= 8'h00;
			14'd2487: ff_rdata <= 8'h00;
			14'd2488: ff_rdata <= 8'h00;
			14'd2489: ff_rdata <= 8'h00;
			14'd2490: ff_rdata <= 8'h00;
			14'd2491: ff_rdata <= 8'h00;
			14'd2492: ff_rdata <= 8'h00;
			14'd2493: ff_rdata <= 8'h00;
			14'd2494: ff_rdata <= 8'h00;
			14'd2495: ff_rdata <= 8'h00;
			14'd2496: ff_rdata <= 8'hFF;
			14'd2497: ff_rdata <= 8'hFF;
			14'd2498: ff_rdata <= 8'hFF;
			14'd2499: ff_rdata <= 8'hFF;
			14'd2500: ff_rdata <= 8'h2C;
			14'd2501: ff_rdata <= 8'hFF;
			14'd2502: ff_rdata <= 8'hFF;
			14'd2503: ff_rdata <= 8'hFF;
			14'd2504: ff_rdata <= 8'hFF;
			14'd2505: ff_rdata <= 8'hFF;
			14'd2506: ff_rdata <= 8'hFF;
			14'd2507: ff_rdata <= 8'hFF;
			14'd2508: ff_rdata <= 8'hFF;
			14'd2509: ff_rdata <= 8'hFF;
			14'd2510: ff_rdata <= 8'hFF;
			14'd2511: ff_rdata <= 8'hFF;
			14'd2512: ff_rdata <= 8'hFF;
			14'd2513: ff_rdata <= 8'hFF;
			14'd2514: ff_rdata <= 8'hFF;
			14'd2515: ff_rdata <= 8'hFF;
			14'd2516: ff_rdata <= 8'hFF;
			14'd2517: ff_rdata <= 8'hFF;
			14'd2518: ff_rdata <= 8'hFF;
			14'd2519: ff_rdata <= 8'hFF;
			14'd2520: ff_rdata <= 8'hFF;
			14'd2521: ff_rdata <= 8'hFF;
			14'd2522: ff_rdata <= 8'hFF;
			14'd2523: ff_rdata <= 8'hFF;
			14'd2524: ff_rdata <= 8'hFF;
			14'd2525: ff_rdata <= 8'h2F;
			14'd2526: ff_rdata <= 8'hFF;
			14'd2527: ff_rdata <= 8'hFF;
			14'd2528: ff_rdata <= 8'hFF;
			14'd2529: ff_rdata <= 8'hFF;
			14'd2530: ff_rdata <= 8'hFF;
			14'd2531: ff_rdata <= 8'hFF;
			14'd2532: ff_rdata <= 8'hFF;
			14'd2533: ff_rdata <= 8'hFF;
			14'd2534: ff_rdata <= 8'hFF;
			14'd2535: ff_rdata <= 8'hFF;
			14'd2536: ff_rdata <= 8'hFF;
			14'd2537: ff_rdata <= 8'hFF;
			14'd2538: ff_rdata <= 8'hFF;
			14'd2539: ff_rdata <= 8'hFF;
			14'd2540: ff_rdata <= 8'hFF;
			14'd2541: ff_rdata <= 8'hFF;
			14'd2542: ff_rdata <= 8'hFF;
			14'd2543: ff_rdata <= 8'hFF;
			14'd2544: ff_rdata <= 8'hFF;
			14'd2545: ff_rdata <= 8'hFF;
			14'd2546: ff_rdata <= 8'hFF;
			14'd2547: ff_rdata <= 8'hFF;
			14'd2548: ff_rdata <= 8'hFF;
			14'd2549: ff_rdata <= 8'hFF;
			14'd2550: ff_rdata <= 8'h32;
			14'd2551: ff_rdata <= 8'hFF;
			14'd2552: ff_rdata <= 8'hFF;
			14'd2553: ff_rdata <= 8'hFF;
			14'd2554: ff_rdata <= 8'hFF;
			14'd2555: ff_rdata <= 8'hFF;
			14'd2556: ff_rdata <= 8'hFF;
			14'd2557: ff_rdata <= 8'hFF;
			14'd2558: ff_rdata <= 8'hFF;
			14'd2559: ff_rdata <= 8'hFF;
			14'd2560: ff_rdata <= 8'h21;
			14'd2561: ff_rdata <= 8'h00;
			14'd2562: ff_rdata <= 8'h00;
			14'd2563: ff_rdata <= 8'h00;
			14'd2564: ff_rdata <= 8'h00;
			14'd2565: ff_rdata <= 8'h00;
			14'd2566: ff_rdata <= 8'h00;
			14'd2567: ff_rdata <= 8'h00;
			14'd2568: ff_rdata <= 8'h00;
			14'd2569: ff_rdata <= 8'h00;
			14'd2570: ff_rdata <= 8'h00;
			14'd2571: ff_rdata <= 8'h00;
			14'd2572: ff_rdata <= 8'h00;
			14'd2573: ff_rdata <= 8'h00;
			14'd2574: ff_rdata <= 8'h00;
			14'd2575: ff_rdata <= 8'h35;
			14'd2576: ff_rdata <= 8'h00;
			14'd2577: ff_rdata <= 8'h00;
			14'd2578: ff_rdata <= 8'h00;
			14'd2579: ff_rdata <= 8'h00;
			14'd2580: ff_rdata <= 8'h00;
			14'd2581: ff_rdata <= 8'h00;
			14'd2582: ff_rdata <= 8'h00;
			14'd2583: ff_rdata <= 8'h00;
			14'd2584: ff_rdata <= 8'h00;
			14'd2585: ff_rdata <= 8'h00;
			14'd2586: ff_rdata <= 8'h00;
			14'd2587: ff_rdata <= 8'h00;
			14'd2588: ff_rdata <= 8'h00;
			14'd2589: ff_rdata <= 8'h00;
			14'd2590: ff_rdata <= 8'h00;
			14'd2591: ff_rdata <= 8'h00;
			14'd2592: ff_rdata <= 8'h00;
			14'd2593: ff_rdata <= 8'h00;
			14'd2594: ff_rdata <= 8'h00;
			14'd2595: ff_rdata <= 8'h00;
			14'd2596: ff_rdata <= 8'h00;
			14'd2597: ff_rdata <= 8'h00;
			14'd2598: ff_rdata <= 8'h00;
			14'd2599: ff_rdata <= 8'h00;
			14'd2600: ff_rdata <= 8'h38;
			14'd2601: ff_rdata <= 8'h00;
			14'd2602: ff_rdata <= 8'h00;
			14'd2603: ff_rdata <= 8'h00;
			14'd2604: ff_rdata <= 8'h00;
			14'd2605: ff_rdata <= 8'h00;
			14'd2606: ff_rdata <= 8'h00;
			14'd2607: ff_rdata <= 8'h00;
			14'd2608: ff_rdata <= 8'h00;
			14'd2609: ff_rdata <= 8'h00;
			14'd2610: ff_rdata <= 8'h00;
			14'd2611: ff_rdata <= 8'h00;
			14'd2612: ff_rdata <= 8'h00;
			14'd2613: ff_rdata <= 8'h00;
			14'd2614: ff_rdata <= 8'h00;
			14'd2615: ff_rdata <= 8'h00;
			14'd2616: ff_rdata <= 8'h00;
			14'd2617: ff_rdata <= 8'h00;
			14'd2618: ff_rdata <= 8'h00;
			14'd2619: ff_rdata <= 8'h00;
			14'd2620: ff_rdata <= 8'h00;
			14'd2621: ff_rdata <= 8'h00;
			14'd2622: ff_rdata <= 8'h00;
			14'd2623: ff_rdata <= 8'h00;
			14'd2624: ff_rdata <= 8'hFF;
			14'd2625: ff_rdata <= 8'h3B;
			14'd2626: ff_rdata <= 8'hFF;
			14'd2627: ff_rdata <= 8'hFF;
			14'd2628: ff_rdata <= 8'hFF;
			14'd2629: ff_rdata <= 8'hFF;
			14'd2630: ff_rdata <= 8'hFF;
			14'd2631: ff_rdata <= 8'hFF;
			14'd2632: ff_rdata <= 8'hFF;
			14'd2633: ff_rdata <= 8'hFF;
			14'd2634: ff_rdata <= 8'hFF;
			14'd2635: ff_rdata <= 8'hFF;
			14'd2636: ff_rdata <= 8'hFF;
			14'd2637: ff_rdata <= 8'hFF;
			14'd2638: ff_rdata <= 8'hFF;
			14'd2639: ff_rdata <= 8'hFF;
			14'd2640: ff_rdata <= 8'hFF;
			14'd2641: ff_rdata <= 8'hFF;
			14'd2642: ff_rdata <= 8'hFF;
			14'd2643: ff_rdata <= 8'hFF;
			14'd2644: ff_rdata <= 8'hFF;
			14'd2645: ff_rdata <= 8'hFF;
			14'd2646: ff_rdata <= 8'hFF;
			14'd2647: ff_rdata <= 8'hFF;
			14'd2648: ff_rdata <= 8'hFF;
			14'd2649: ff_rdata <= 8'hFF;
			14'd2650: ff_rdata <= 8'h3E;
			14'd2651: ff_rdata <= 8'hFF;
			14'd2652: ff_rdata <= 8'hFF;
			14'd2653: ff_rdata <= 8'hFF;
			14'd2654: ff_rdata <= 8'hFF;
			14'd2655: ff_rdata <= 8'hFF;
			14'd2656: ff_rdata <= 8'hFF;
			14'd2657: ff_rdata <= 8'hFF;
			14'd2658: ff_rdata <= 8'hFF;
			14'd2659: ff_rdata <= 8'hFF;
			14'd2660: ff_rdata <= 8'hFF;
			14'd2661: ff_rdata <= 8'hFF;
			14'd2662: ff_rdata <= 8'hFF;
			14'd2663: ff_rdata <= 8'hFF;
			14'd2664: ff_rdata <= 8'hFF;
			14'd2665: ff_rdata <= 8'hFF;
			14'd2666: ff_rdata <= 8'hFF;
			14'd2667: ff_rdata <= 8'hFF;
			14'd2668: ff_rdata <= 8'hFF;
			14'd2669: ff_rdata <= 8'hFF;
			14'd2670: ff_rdata <= 8'hFF;
			14'd2671: ff_rdata <= 8'hFF;
			14'd2672: ff_rdata <= 8'hFF;
			14'd2673: ff_rdata <= 8'hFF;
			14'd2674: ff_rdata <= 8'hFF;
			14'd2675: ff_rdata <= 8'h41;
			14'd2676: ff_rdata <= 8'hFF;
			14'd2677: ff_rdata <= 8'hFF;
			14'd2678: ff_rdata <= 8'hFF;
			14'd2679: ff_rdata <= 8'hFF;
			14'd2680: ff_rdata <= 8'hFF;
			14'd2681: ff_rdata <= 8'hFF;
			14'd2682: ff_rdata <= 8'hFF;
			14'd2683: ff_rdata <= 8'hFF;
			14'd2684: ff_rdata <= 8'hFF;
			14'd2685: ff_rdata <= 8'hFF;
			14'd2686: ff_rdata <= 8'hFF;
			14'd2687: ff_rdata <= 8'h3F;
			14'd2688: ff_rdata <= 8'h01;
			14'd2689: ff_rdata <= 8'h00;
			14'd2690: ff_rdata <= 8'h00;
			14'd2691: ff_rdata <= 8'h00;
			14'd2692: ff_rdata <= 8'h00;
			14'd2693: ff_rdata <= 8'h00;
			14'd2694: ff_rdata <= 8'h00;
			14'd2695: ff_rdata <= 8'h00;
			14'd2696: ff_rdata <= 8'h00;
			14'd2697: ff_rdata <= 8'h00;
			14'd2698: ff_rdata <= 8'h00;
			14'd2699: ff_rdata <= 8'h00;
			14'd2700: ff_rdata <= 8'h44;
			14'd2701: ff_rdata <= 8'h00;
			14'd2702: ff_rdata <= 8'h00;
			14'd2703: ff_rdata <= 8'h00;
			14'd2704: ff_rdata <= 8'h00;
			14'd2705: ff_rdata <= 8'h00;
			14'd2706: ff_rdata <= 8'h00;
			14'd2707: ff_rdata <= 8'h00;
			14'd2708: ff_rdata <= 8'h00;
			14'd2709: ff_rdata <= 8'h00;
			14'd2710: ff_rdata <= 8'h00;
			14'd2711: ff_rdata <= 8'h00;
			14'd2712: ff_rdata <= 8'h00;
			14'd2713: ff_rdata <= 8'h00;
			14'd2714: ff_rdata <= 8'h00;
			14'd2715: ff_rdata <= 8'h00;
			14'd2716: ff_rdata <= 8'h00;
			14'd2717: ff_rdata <= 8'h00;
			14'd2718: ff_rdata <= 8'h00;
			14'd2719: ff_rdata <= 8'h00;
			14'd2720: ff_rdata <= 8'h00;
			14'd2721: ff_rdata <= 8'h00;
			14'd2722: ff_rdata <= 8'h00;
			14'd2723: ff_rdata <= 8'h00;
			14'd2724: ff_rdata <= 8'h00;
			14'd2725: ff_rdata <= 8'h47;
			14'd2726: ff_rdata <= 8'h00;
			14'd2727: ff_rdata <= 8'h00;
			14'd2728: ff_rdata <= 8'h00;
			14'd2729: ff_rdata <= 8'h00;
			14'd2730: ff_rdata <= 8'h00;
			14'd2731: ff_rdata <= 8'h00;
			14'd2732: ff_rdata <= 8'h00;
			14'd2733: ff_rdata <= 8'h00;
			14'd2734: ff_rdata <= 8'h00;
			14'd2735: ff_rdata <= 8'h00;
			14'd2736: ff_rdata <= 8'h00;
			14'd2737: ff_rdata <= 8'h00;
			14'd2738: ff_rdata <= 8'h00;
			14'd2739: ff_rdata <= 8'h00;
			14'd2740: ff_rdata <= 8'h00;
			14'd2741: ff_rdata <= 8'h00;
			14'd2742: ff_rdata <= 8'h00;
			14'd2743: ff_rdata <= 8'h00;
			14'd2744: ff_rdata <= 8'h00;
			14'd2745: ff_rdata <= 8'h00;
			14'd2746: ff_rdata <= 8'h00;
			14'd2747: ff_rdata <= 8'h00;
			14'd2748: ff_rdata <= 8'h00;
			14'd2749: ff_rdata <= 8'h00;
			14'd2750: ff_rdata <= 8'h4A;
			14'd2751: ff_rdata <= 8'h00;
			14'd2752: ff_rdata <= 8'hFF;
			14'd2753: ff_rdata <= 8'hFF;
			14'd2754: ff_rdata <= 8'hFF;
			14'd2755: ff_rdata <= 8'hFF;
			14'd2756: ff_rdata <= 8'hFF;
			14'd2757: ff_rdata <= 8'hFF;
			14'd2758: ff_rdata <= 8'hFF;
			14'd2759: ff_rdata <= 8'hFF;
			14'd2760: ff_rdata <= 8'hFF;
			14'd2761: ff_rdata <= 8'hFF;
			14'd2762: ff_rdata <= 8'hFF;
			14'd2763: ff_rdata <= 8'hFF;
			14'd2764: ff_rdata <= 8'hFF;
			14'd2765: ff_rdata <= 8'hFF;
			14'd2766: ff_rdata <= 8'hFF;
			14'd2767: ff_rdata <= 8'hFF;
			14'd2768: ff_rdata <= 8'hFF;
			14'd2769: ff_rdata <= 8'hFF;
			14'd2770: ff_rdata <= 8'hFF;
			14'd2771: ff_rdata <= 8'hFF;
			14'd2772: ff_rdata <= 8'hFF;
			14'd2773: ff_rdata <= 8'hFF;
			14'd2774: ff_rdata <= 8'hFF;
			14'd2775: ff_rdata <= 8'h4D;
			14'd2776: ff_rdata <= 8'hFF;
			14'd2777: ff_rdata <= 8'hFF;
			14'd2778: ff_rdata <= 8'hFF;
			14'd2779: ff_rdata <= 8'hFF;
			14'd2780: ff_rdata <= 8'hFF;
			14'd2781: ff_rdata <= 8'hFF;
			14'd2782: ff_rdata <= 8'hFF;
			14'd2783: ff_rdata <= 8'hFF;
			14'd2784: ff_rdata <= 8'hFF;
			14'd2785: ff_rdata <= 8'hFF;
			14'd2786: ff_rdata <= 8'hFF;
			14'd2787: ff_rdata <= 8'hFF;
			14'd2788: ff_rdata <= 8'hFF;
			14'd2789: ff_rdata <= 8'hFF;
			14'd2790: ff_rdata <= 8'hFF;
			14'd2791: ff_rdata <= 8'hFF;
			14'd2792: ff_rdata <= 8'hFF;
			14'd2793: ff_rdata <= 8'hFF;
			14'd2794: ff_rdata <= 8'hFF;
			14'd2795: ff_rdata <= 8'hFF;
			14'd2796: ff_rdata <= 8'hFF;
			14'd2797: ff_rdata <= 8'hFF;
			14'd2798: ff_rdata <= 8'hFF;
			14'd2799: ff_rdata <= 8'hFF;
			14'd2800: ff_rdata <= 8'h50;
			14'd2801: ff_rdata <= 8'hFF;
			14'd2802: ff_rdata <= 8'hFF;
			14'd2803: ff_rdata <= 8'hFF;
			14'd2804: ff_rdata <= 8'hFF;
			14'd2805: ff_rdata <= 8'hFF;
			14'd2806: ff_rdata <= 8'hFF;
			14'd2807: ff_rdata <= 8'hFF;
			14'd2808: ff_rdata <= 8'hFF;
			14'd2809: ff_rdata <= 8'hFF;
			14'd2810: ff_rdata <= 8'hFF;
			14'd2811: ff_rdata <= 8'hFF;
			14'd2812: ff_rdata <= 8'hFF;
			14'd2813: ff_rdata <= 8'hFF;
			14'd2814: ff_rdata <= 8'hFF;
			14'd2815: ff_rdata <= 8'hFF;
			14'd2816: ff_rdata <= 8'hFF;
			14'd2817: ff_rdata <= 8'hFF;
			14'd2818: ff_rdata <= 8'hFF;
			14'd2819: ff_rdata <= 8'hFF;
			14'd2820: ff_rdata <= 8'hFF;
			14'd2821: ff_rdata <= 8'hFF;
			14'd2822: ff_rdata <= 8'hFF;
			14'd2823: ff_rdata <= 8'hFF;
			14'd2824: ff_rdata <= 8'hFF;
			14'd2825: ff_rdata <= 8'h53;
			14'd2826: ff_rdata <= 8'hFF;
			14'd2827: ff_rdata <= 8'hFF;
			14'd2828: ff_rdata <= 8'hFF;
			14'd2829: ff_rdata <= 8'hFF;
			14'd2830: ff_rdata <= 8'hFF;
			14'd2831: ff_rdata <= 8'hFF;
			14'd2832: ff_rdata <= 8'hFF;
			14'd2833: ff_rdata <= 8'hFF;
			14'd2834: ff_rdata <= 8'hFF;
			14'd2835: ff_rdata <= 8'hFF;
			14'd2836: ff_rdata <= 8'hFF;
			14'd2837: ff_rdata <= 8'hFF;
			14'd2838: ff_rdata <= 8'hFF;
			14'd2839: ff_rdata <= 8'hFF;
			14'd2840: ff_rdata <= 8'hFF;
			14'd2841: ff_rdata <= 8'hFF;
			14'd2842: ff_rdata <= 8'hFF;
			14'd2843: ff_rdata <= 8'hFF;
			14'd2844: ff_rdata <= 8'hFF;
			14'd2845: ff_rdata <= 8'hFF;
			14'd2846: ff_rdata <= 8'hFF;
			14'd2847: ff_rdata <= 8'hFF;
			14'd2848: ff_rdata <= 8'hFF;
			14'd2849: ff_rdata <= 8'hFF;
			14'd2850: ff_rdata <= 8'h56;
			14'd2851: ff_rdata <= 8'hFF;
			14'd2852: ff_rdata <= 8'hFF;
			14'd2853: ff_rdata <= 8'hFF;
			14'd2854: ff_rdata <= 8'hFF;
			14'd2855: ff_rdata <= 8'hFF;
			14'd2856: ff_rdata <= 8'hFF;
			14'd2857: ff_rdata <= 8'hFF;
			14'd2858: ff_rdata <= 8'hFF;
			14'd2859: ff_rdata <= 8'hFF;
			14'd2860: ff_rdata <= 8'hFF;
			14'd2861: ff_rdata <= 8'hFF;
			14'd2862: ff_rdata <= 8'hFF;
			14'd2863: ff_rdata <= 8'hFF;
			14'd2864: ff_rdata <= 8'hFF;
			14'd2865: ff_rdata <= 8'hFF;
			14'd2866: ff_rdata <= 8'hFF;
			14'd2867: ff_rdata <= 8'hFF;
			14'd2868: ff_rdata <= 8'hFF;
			14'd2869: ff_rdata <= 8'hFF;
			14'd2870: ff_rdata <= 8'hFF;
			14'd2871: ff_rdata <= 8'hFF;
			14'd2872: ff_rdata <= 8'hFF;
			14'd2873: ff_rdata <= 8'hFF;
			14'd2874: ff_rdata <= 8'hFF;
			14'd2875: ff_rdata <= 8'h59;
			14'd2876: ff_rdata <= 8'hFF;
			14'd2877: ff_rdata <= 8'hFF;
			14'd2878: ff_rdata <= 8'hFF;
			14'd2879: ff_rdata <= 8'hFF;
			14'd2880: ff_rdata <= 8'h00;
			14'd2881: ff_rdata <= 8'h00;
			14'd2882: ff_rdata <= 8'h00;
			14'd2883: ff_rdata <= 8'h00;
			14'd2884: ff_rdata <= 8'h00;
			14'd2885: ff_rdata <= 8'h00;
			14'd2886: ff_rdata <= 8'h00;
			14'd2887: ff_rdata <= 8'h00;
			14'd2888: ff_rdata <= 8'h00;
			14'd2889: ff_rdata <= 8'h00;
			14'd2890: ff_rdata <= 8'h00;
			14'd2891: ff_rdata <= 8'h00;
			14'd2892: ff_rdata <= 8'h00;
			14'd2893: ff_rdata <= 8'h00;
			14'd2894: ff_rdata <= 8'h00;
			14'd2895: ff_rdata <= 8'h00;
			14'd2896: ff_rdata <= 8'h00;
			14'd2897: ff_rdata <= 8'h00;
			14'd2898: ff_rdata <= 8'h00;
			14'd2899: ff_rdata <= 8'h00;
			14'd2900: ff_rdata <= 8'h5C;
			14'd2901: ff_rdata <= 8'h00;
			14'd2902: ff_rdata <= 8'h00;
			14'd2903: ff_rdata <= 8'h00;
			14'd2904: ff_rdata <= 8'h00;
			14'd2905: ff_rdata <= 8'h00;
			14'd2906: ff_rdata <= 8'h00;
			14'd2907: ff_rdata <= 8'h00;
			14'd2908: ff_rdata <= 8'h00;
			14'd2909: ff_rdata <= 8'h00;
			14'd2910: ff_rdata <= 8'h00;
			14'd2911: ff_rdata <= 8'h00;
			14'd2912: ff_rdata <= 8'h00;
			14'd2913: ff_rdata <= 8'h00;
			14'd2914: ff_rdata <= 8'h00;
			14'd2915: ff_rdata <= 8'h00;
			14'd2916: ff_rdata <= 8'h00;
			14'd2917: ff_rdata <= 8'h00;
			14'd2918: ff_rdata <= 8'h00;
			14'd2919: ff_rdata <= 8'h00;
			14'd2920: ff_rdata <= 8'h00;
			14'd2921: ff_rdata <= 8'h00;
			14'd2922: ff_rdata <= 8'h00;
			14'd2923: ff_rdata <= 8'h00;
			14'd2924: ff_rdata <= 8'h00;
			14'd2925: ff_rdata <= 8'h5F;
			14'd2926: ff_rdata <= 8'h00;
			14'd2927: ff_rdata <= 8'h00;
			14'd2928: ff_rdata <= 8'h00;
			14'd2929: ff_rdata <= 8'h00;
			14'd2930: ff_rdata <= 8'h00;
			14'd2931: ff_rdata <= 8'h00;
			14'd2932: ff_rdata <= 8'h00;
			14'd2933: ff_rdata <= 8'h00;
			14'd2934: ff_rdata <= 8'h00;
			14'd2935: ff_rdata <= 8'h00;
			14'd2936: ff_rdata <= 8'h00;
			14'd2937: ff_rdata <= 8'h00;
			14'd2938: ff_rdata <= 8'h00;
			14'd2939: ff_rdata <= 8'h00;
			14'd2940: ff_rdata <= 8'h00;
			14'd2941: ff_rdata <= 8'h00;
			14'd2942: ff_rdata <= 8'h00;
			14'd2943: ff_rdata <= 8'h89;
			14'd2944: ff_rdata <= 8'hDF;
			14'd2945: ff_rdata <= 8'hFF;
			14'd2946: ff_rdata <= 8'hFF;
			14'd2947: ff_rdata <= 8'hFF;
			14'd2948: ff_rdata <= 8'hFF;
			14'd2949: ff_rdata <= 8'hFF;
			14'd2950: ff_rdata <= 8'h62;
			14'd2951: ff_rdata <= 8'hFF;
			14'd2952: ff_rdata <= 8'hFF;
			14'd2953: ff_rdata <= 8'hFF;
			14'd2954: ff_rdata <= 8'hFF;
			14'd2955: ff_rdata <= 8'hFF;
			14'd2956: ff_rdata <= 8'hFF;
			14'd2957: ff_rdata <= 8'hFF;
			14'd2958: ff_rdata <= 8'hFF;
			14'd2959: ff_rdata <= 8'hFF;
			14'd2960: ff_rdata <= 8'hFF;
			14'd2961: ff_rdata <= 8'hFF;
			14'd2962: ff_rdata <= 8'hFF;
			14'd2963: ff_rdata <= 8'hFF;
			14'd2964: ff_rdata <= 8'hFF;
			14'd2965: ff_rdata <= 8'hFF;
			14'd2966: ff_rdata <= 8'hFF;
			14'd2967: ff_rdata <= 8'hFF;
			14'd2968: ff_rdata <= 8'hFF;
			14'd2969: ff_rdata <= 8'hFF;
			14'd2970: ff_rdata <= 8'hFF;
			14'd2971: ff_rdata <= 8'hFF;
			14'd2972: ff_rdata <= 8'hFF;
			14'd2973: ff_rdata <= 8'hFF;
			14'd2974: ff_rdata <= 8'hFF;
			14'd2975: ff_rdata <= 8'h65;
			14'd2976: ff_rdata <= 8'hFF;
			14'd2977: ff_rdata <= 8'hFF;
			14'd2978: ff_rdata <= 8'hFF;
			14'd2979: ff_rdata <= 8'hFF;
			14'd2980: ff_rdata <= 8'hFF;
			14'd2981: ff_rdata <= 8'hFF;
			14'd2982: ff_rdata <= 8'hFF;
			14'd2983: ff_rdata <= 8'hFF;
			14'd2984: ff_rdata <= 8'hFF;
			14'd2985: ff_rdata <= 8'hFF;
			14'd2986: ff_rdata <= 8'hFF;
			14'd2987: ff_rdata <= 8'hFF;
			14'd2988: ff_rdata <= 8'hFF;
			14'd2989: ff_rdata <= 8'hFF;
			14'd2990: ff_rdata <= 8'hFF;
			14'd2991: ff_rdata <= 8'hFF;
			14'd2992: ff_rdata <= 8'hFF;
			14'd2993: ff_rdata <= 8'hFF;
			14'd2994: ff_rdata <= 8'hFF;
			14'd2995: ff_rdata <= 8'hFF;
			14'd2996: ff_rdata <= 8'hFF;
			14'd2997: ff_rdata <= 8'hFF;
			14'd2998: ff_rdata <= 8'hFF;
			14'd2999: ff_rdata <= 8'hFF;
			14'd3000: ff_rdata <= 8'h68;
			14'd3001: ff_rdata <= 8'hFF;
			14'd3002: ff_rdata <= 8'hFF;
			14'd3003: ff_rdata <= 8'hFF;
			14'd3004: ff_rdata <= 8'hFF;
			14'd3005: ff_rdata <= 8'hFF;
			14'd3006: ff_rdata <= 8'hFF;
			14'd3007: ff_rdata <= 8'hFF;
			14'd3008: ff_rdata <= 8'h00;
			14'd3009: ff_rdata <= 8'h00;
			14'd3010: ff_rdata <= 8'h00;
			14'd3011: ff_rdata <= 8'h00;
			14'd3012: ff_rdata <= 8'h00;
			14'd3013: ff_rdata <= 8'h00;
			14'd3014: ff_rdata <= 8'h00;
			14'd3015: ff_rdata <= 8'h00;
			14'd3016: ff_rdata <= 8'h00;
			14'd3017: ff_rdata <= 8'h00;
			14'd3018: ff_rdata <= 8'h00;
			14'd3019: ff_rdata <= 8'h00;
			14'd3020: ff_rdata <= 8'h00;
			14'd3021: ff_rdata <= 8'h00;
			14'd3022: ff_rdata <= 8'h00;
			14'd3023: ff_rdata <= 8'h00;
			14'd3024: ff_rdata <= 8'h00;
			14'd3025: ff_rdata <= 8'h6B;
			14'd3026: ff_rdata <= 8'h00;
			14'd3027: ff_rdata <= 8'h00;
			14'd3028: ff_rdata <= 8'h00;
			14'd3029: ff_rdata <= 8'h00;
			14'd3030: ff_rdata <= 8'h00;
			14'd3031: ff_rdata <= 8'h00;
			14'd3032: ff_rdata <= 8'h00;
			14'd3033: ff_rdata <= 8'h00;
			14'd3034: ff_rdata <= 8'h00;
			14'd3035: ff_rdata <= 8'h00;
			14'd3036: ff_rdata <= 8'h00;
			14'd3037: ff_rdata <= 8'h00;
			14'd3038: ff_rdata <= 8'h00;
			14'd3039: ff_rdata <= 8'h00;
			14'd3040: ff_rdata <= 8'h00;
			14'd3041: ff_rdata <= 8'h00;
			14'd3042: ff_rdata <= 8'h00;
			14'd3043: ff_rdata <= 8'h00;
			14'd3044: ff_rdata <= 8'h00;
			14'd3045: ff_rdata <= 8'h00;
			14'd3046: ff_rdata <= 8'h00;
			14'd3047: ff_rdata <= 8'h00;
			14'd3048: ff_rdata <= 8'h00;
			14'd3049: ff_rdata <= 8'h00;
			14'd3050: ff_rdata <= 8'h6E;
			14'd3051: ff_rdata <= 8'h00;
			14'd3052: ff_rdata <= 8'h00;
			14'd3053: ff_rdata <= 8'h00;
			14'd3054: ff_rdata <= 8'h00;
			14'd3055: ff_rdata <= 8'h00;
			14'd3056: ff_rdata <= 8'h00;
			14'd3057: ff_rdata <= 8'h00;
			14'd3058: ff_rdata <= 8'h00;
			14'd3059: ff_rdata <= 8'h00;
			14'd3060: ff_rdata <= 8'h00;
			14'd3061: ff_rdata <= 8'h00;
			14'd3062: ff_rdata <= 8'h00;
			14'd3063: ff_rdata <= 8'h00;
			14'd3064: ff_rdata <= 8'h00;
			14'd3065: ff_rdata <= 8'h00;
			14'd3066: ff_rdata <= 8'h00;
			14'd3067: ff_rdata <= 8'h00;
			14'd3068: ff_rdata <= 8'h00;
			14'd3069: ff_rdata <= 8'h00;
			14'd3070: ff_rdata <= 8'h00;
			14'd3071: ff_rdata <= 8'h00;
			14'd3072: ff_rdata <= 8'h31;
			14'd3073: ff_rdata <= 8'h11;
			14'd3074: ff_rdata <= 8'h0E;
			14'd3075: ff_rdata <= 8'h20;
			14'd3076: ff_rdata <= 8'hD9;
			14'd3077: ff_rdata <= 8'hB2;
			14'd3078: ff_rdata <= 8'h11;
			14'd3079: ff_rdata <= 8'hF4;
			14'd3080: ff_rdata <= 8'h30;
			14'd3081: ff_rdata <= 8'h10;
			14'd3082: ff_rdata <= 8'h0F;
			14'd3083: ff_rdata <= 8'h20;
			14'd3084: ff_rdata <= 8'hD9;
			14'd3085: ff_rdata <= 8'hB2;
			14'd3086: ff_rdata <= 8'h10;
			14'd3087: ff_rdata <= 8'hF3;
			14'd3088: ff_rdata <= 8'h61;
			14'd3089: ff_rdata <= 8'h61;
			14'd3090: ff_rdata <= 8'h12;
			14'd3091: ff_rdata <= 8'h20;
			14'd3092: ff_rdata <= 8'hB4;
			14'd3093: ff_rdata <= 8'h56;
			14'd3094: ff_rdata <= 8'h14;
			14'd3095: ff_rdata <= 8'h17;
			14'd3096: ff_rdata <= 8'h61;
			14'd3097: ff_rdata <= 8'h31;
			14'd3098: ff_rdata <= 8'h20;
			14'd3099: ff_rdata <= 8'h20;
			14'd3100: ff_rdata <= 8'h6C;
			14'd3101: ff_rdata <= 8'h43;
			14'd3102: ff_rdata <= 8'h18;
			14'd3103: ff_rdata <= 8'h26;
			14'd3104: ff_rdata <= 8'hA2;
			14'd3105: ff_rdata <= 8'h30;
			14'd3106: ff_rdata <= 8'hA0;
			14'd3107: ff_rdata <= 8'h20;
			14'd3108: ff_rdata <= 8'h88;
			14'd3109: ff_rdata <= 8'h54;
			14'd3110: ff_rdata <= 8'h14;
			14'd3111: ff_rdata <= 8'h06;
			14'd3112: ff_rdata <= 8'h31;
			14'd3113: ff_rdata <= 8'h34;
			14'd3114: ff_rdata <= 8'h20;
			14'd3115: ff_rdata <= 8'h20;
			14'd3116: ff_rdata <= 8'h72;
			14'd3117: ff_rdata <= 8'h56;
			14'd3118: ff_rdata <= 8'h0A;
			14'd3119: ff_rdata <= 8'h1C;
			14'd3120: ff_rdata <= 8'h31;
			14'd3121: ff_rdata <= 8'h71;
			14'd3122: ff_rdata <= 8'h16;
			14'd3123: ff_rdata <= 8'h20;
			14'd3124: ff_rdata <= 8'h51;
			14'd3125: ff_rdata <= 8'h52;
			14'd3126: ff_rdata <= 8'h26;
			14'd3127: ff_rdata <= 8'h24;
			14'd3128: ff_rdata <= 8'h34;
			14'd3129: ff_rdata <= 8'h30;
			14'd3130: ff_rdata <= 8'h37;
			14'd3131: ff_rdata <= 8'h20;
			14'd3132: ff_rdata <= 8'h50;
			14'd3133: ff_rdata <= 8'h30;
			14'd3134: ff_rdata <= 8'h76;
			14'd3135: ff_rdata <= 8'h06;
			14'd3136: ff_rdata <= 8'h17;
			14'd3137: ff_rdata <= 8'h52;
			14'd3138: ff_rdata <= 8'h18;
			14'd3139: ff_rdata <= 8'h20;
			14'd3140: ff_rdata <= 8'h88;
			14'd3141: ff_rdata <= 8'hD9;
			14'd3142: ff_rdata <= 8'h66;
			14'd3143: ff_rdata <= 8'h24;
			14'd3144: ff_rdata <= 8'hE1;
			14'd3145: ff_rdata <= 8'h63;
			14'd3146: ff_rdata <= 8'h0A;
			14'd3147: ff_rdata <= 8'h20;
			14'd3148: ff_rdata <= 8'hFC;
			14'd3149: ff_rdata <= 8'hF8;
			14'd3150: ff_rdata <= 8'h28;
			14'd3151: ff_rdata <= 8'h29;
			14'd3152: ff_rdata <= 8'h02;
			14'd3153: ff_rdata <= 8'h41;
			14'd3154: ff_rdata <= 8'h15;
			14'd3155: ff_rdata <= 8'h20;
			14'd3156: ff_rdata <= 8'hA3;
			14'd3157: ff_rdata <= 8'hA3;
			14'd3158: ff_rdata <= 8'h75;
			14'd3159: ff_rdata <= 8'h05;
			14'd3160: ff_rdata <= 8'h19;
			14'd3161: ff_rdata <= 8'h53;
			14'd3162: ff_rdata <= 8'h0C;
			14'd3163: ff_rdata <= 8'h20;
			14'd3164: ff_rdata <= 8'hC7;
			14'd3165: ff_rdata <= 8'hF5;
			14'd3166: ff_rdata <= 8'h11;
			14'd3167: ff_rdata <= 8'h03;
			14'd3168: ff_rdata <= 8'h23;
			14'd3169: ff_rdata <= 8'h43;
			14'd3170: ff_rdata <= 8'h09;
			14'd3171: ff_rdata <= 8'h20;
			14'd3172: ff_rdata <= 8'hDD;
			14'd3173: ff_rdata <= 8'hBF;
			14'd3174: ff_rdata <= 8'h4A;
			14'd3175: ff_rdata <= 8'h05;
			14'd3176: ff_rdata <= 8'h03;
			14'd3177: ff_rdata <= 8'h09;
			14'd3178: ff_rdata <= 8'h11;
			14'd3179: ff_rdata <= 8'h20;
			14'd3180: ff_rdata <= 8'hD2;
			14'd3181: ff_rdata <= 8'hB4;
			14'd3182: ff_rdata <= 8'hF4;
			14'd3183: ff_rdata <= 8'hF5;
			14'd3184: ff_rdata <= 8'h01;
			14'd3185: ff_rdata <= 8'h00;
			14'd3186: ff_rdata <= 8'h06;
			14'd3187: ff_rdata <= 8'h20;
			14'd3188: ff_rdata <= 8'hA3;
			14'd3189: ff_rdata <= 8'hE2;
			14'd3190: ff_rdata <= 8'hF4;
			14'd3191: ff_rdata <= 8'hF4;
			14'd3192: ff_rdata <= 8'h01;
			14'd3193: ff_rdata <= 8'h01;
			14'd3194: ff_rdata <= 8'h11;
			14'd3195: ff_rdata <= 8'h20;
			14'd3196: ff_rdata <= 8'hC0;
			14'd3197: ff_rdata <= 8'hB4;
			14'd3198: ff_rdata <= 8'h01;
			14'd3199: ff_rdata <= 8'hF6;
			14'd3200: ff_rdata <= 8'hF9;
			14'd3201: ff_rdata <= 8'hF1;
			14'd3202: ff_rdata <= 8'h24;
			14'd3203: ff_rdata <= 8'h20;
			14'd3204: ff_rdata <= 8'h95;
			14'd3205: ff_rdata <= 8'hD1;
			14'd3206: ff_rdata <= 8'hE5;
			14'd3207: ff_rdata <= 8'hF2;
			14'd3208: ff_rdata <= 8'h13;
			14'd3209: ff_rdata <= 8'h11;
			14'd3210: ff_rdata <= 8'h0C;
			14'd3211: ff_rdata <= 8'h20;
			14'd3212: ff_rdata <= 8'hFC;
			14'd3213: ff_rdata <= 8'hD2;
			14'd3214: ff_rdata <= 8'h33;
			14'd3215: ff_rdata <= 8'h83;
			14'd3216: ff_rdata <= 8'h01;
			14'd3217: ff_rdata <= 8'h10;
			14'd3218: ff_rdata <= 8'h0E;
			14'd3219: ff_rdata <= 8'h20;
			14'd3220: ff_rdata <= 8'hCA;
			14'd3221: ff_rdata <= 8'hE6;
			14'd3222: ff_rdata <= 8'h44;
			14'd3223: ff_rdata <= 8'h24;
			14'd3224: ff_rdata <= 8'hE0;
			14'd3225: ff_rdata <= 8'hF4;
			14'd3226: ff_rdata <= 8'h1B;
			14'd3227: ff_rdata <= 8'h20;
			14'd3228: ff_rdata <= 8'h11;
			14'd3229: ff_rdata <= 8'hF0;
			14'd3230: ff_rdata <= 8'h04;
			14'd3231: ff_rdata <= 8'h08;
			14'd3232: ff_rdata <= 8'hFF;
			14'd3233: ff_rdata <= 8'h70;
			14'd3234: ff_rdata <= 8'h19;
			14'd3235: ff_rdata <= 8'h20;
			14'd3236: ff_rdata <= 8'h50;
			14'd3237: ff_rdata <= 8'h1F;
			14'd3238: ff_rdata <= 8'h05;
			14'd3239: ff_rdata <= 8'h01;
			14'd3240: ff_rdata <= 8'h13;
			14'd3241: ff_rdata <= 8'h11;
			14'd3242: ff_rdata <= 8'h11;
			14'd3243: ff_rdata <= 8'h20;
			14'd3244: ff_rdata <= 8'hFA;
			14'd3245: ff_rdata <= 8'hF2;
			14'd3246: ff_rdata <= 8'h21;
			14'd3247: ff_rdata <= 8'hF4;
			14'd3248: ff_rdata <= 8'hA6;
			14'd3249: ff_rdata <= 8'h42;
			14'd3250: ff_rdata <= 8'h10;
			14'd3251: ff_rdata <= 8'h20;
			14'd3252: ff_rdata <= 8'hFB;
			14'd3253: ff_rdata <= 8'hB9;
			14'd3254: ff_rdata <= 8'h11;
			14'd3255: ff_rdata <= 8'h02;
			14'd3256: ff_rdata <= 8'h40;
			14'd3257: ff_rdata <= 8'h31;
			14'd3258: ff_rdata <= 8'h89;
			14'd3259: ff_rdata <= 8'h20;
			14'd3260: ff_rdata <= 8'hC7;
			14'd3261: ff_rdata <= 8'hF9;
			14'd3262: ff_rdata <= 8'h14;
			14'd3263: ff_rdata <= 8'h04;
			14'd3264: ff_rdata <= 8'h42;
			14'd3265: ff_rdata <= 8'h44;
			14'd3266: ff_rdata <= 8'h0B;
			14'd3267: ff_rdata <= 8'h20;
			14'd3268: ff_rdata <= 8'h94;
			14'd3269: ff_rdata <= 8'hB0;
			14'd3270: ff_rdata <= 8'h33;
			14'd3271: ff_rdata <= 8'hF6;
			14'd3272: ff_rdata <= 8'h01;
			14'd3273: ff_rdata <= 8'h03;
			14'd3274: ff_rdata <= 8'h0B;
			14'd3275: ff_rdata <= 8'h20;
			14'd3276: ff_rdata <= 8'hBA;
			14'd3277: ff_rdata <= 8'hD9;
			14'd3278: ff_rdata <= 8'h25;
			14'd3279: ff_rdata <= 8'h06;
			14'd3280: ff_rdata <= 8'h40;
			14'd3281: ff_rdata <= 8'h00;
			14'd3282: ff_rdata <= 8'h00;
			14'd3283: ff_rdata <= 8'h20;
			14'd3284: ff_rdata <= 8'hFA;
			14'd3285: ff_rdata <= 8'hD9;
			14'd3286: ff_rdata <= 8'h37;
			14'd3287: ff_rdata <= 8'h04;
			14'd3288: ff_rdata <= 8'h02;
			14'd3289: ff_rdata <= 8'h03;
			14'd3290: ff_rdata <= 8'h09;
			14'd3291: ff_rdata <= 8'h20;
			14'd3292: ff_rdata <= 8'hCB;
			14'd3293: ff_rdata <= 8'hFF;
			14'd3294: ff_rdata <= 8'h39;
			14'd3295: ff_rdata <= 8'h06;
			14'd3296: ff_rdata <= 8'h18;
			14'd3297: ff_rdata <= 8'h11;
			14'd3298: ff_rdata <= 8'h09;
			14'd3299: ff_rdata <= 8'h20;
			14'd3300: ff_rdata <= 8'hF8;
			14'd3301: ff_rdata <= 8'hF5;
			14'd3302: ff_rdata <= 8'h26;
			14'd3303: ff_rdata <= 8'h26;
			14'd3304: ff_rdata <= 8'h0B;
			14'd3305: ff_rdata <= 8'h04;
			14'd3306: ff_rdata <= 8'h09;
			14'd3307: ff_rdata <= 8'h20;
			14'd3308: ff_rdata <= 8'hF0;
			14'd3309: ff_rdata <= 8'hF5;
			14'd3310: ff_rdata <= 8'h01;
			14'd3311: ff_rdata <= 8'h27;
			14'd3312: ff_rdata <= 8'h40;
			14'd3313: ff_rdata <= 8'h40;
			14'd3314: ff_rdata <= 8'h07;
			14'd3315: ff_rdata <= 8'h20;
			14'd3316: ff_rdata <= 8'hD0;
			14'd3317: ff_rdata <= 8'hD6;
			14'd3318: ff_rdata <= 8'h01;
			14'd3319: ff_rdata <= 8'h27;
			14'd3320: ff_rdata <= 8'h00;
			14'd3321: ff_rdata <= 8'h01;
			14'd3322: ff_rdata <= 8'h07;
			14'd3323: ff_rdata <= 8'h20;
			14'd3324: ff_rdata <= 8'hCB;
			14'd3325: ff_rdata <= 8'hE3;
			14'd3326: ff_rdata <= 8'h36;
			14'd3327: ff_rdata <= 8'h25;
			14'd3328: ff_rdata <= 8'h11;
			14'd3329: ff_rdata <= 8'h11;
			14'd3330: ff_rdata <= 8'h08;
			14'd3331: ff_rdata <= 8'h20;
			14'd3332: ff_rdata <= 8'hFA;
			14'd3333: ff_rdata <= 8'hB2;
			14'd3334: ff_rdata <= 8'h20;
			14'd3335: ff_rdata <= 8'hF4;
			14'd3336: ff_rdata <= 8'h11;
			14'd3337: ff_rdata <= 8'h11;
			14'd3338: ff_rdata <= 8'h11;
			14'd3339: ff_rdata <= 8'h20;
			14'd3340: ff_rdata <= 8'hC0;
			14'd3341: ff_rdata <= 8'hB2;
			14'd3342: ff_rdata <= 8'h01;
			14'd3343: ff_rdata <= 8'hF4;
			14'd3344: ff_rdata <= 8'h19;
			14'd3345: ff_rdata <= 8'h53;
			14'd3346: ff_rdata <= 8'h15;
			14'd3347: ff_rdata <= 8'h20;
			14'd3348: ff_rdata <= 8'hE7;
			14'd3349: ff_rdata <= 8'h95;
			14'd3350: ff_rdata <= 8'h21;
			14'd3351: ff_rdata <= 8'h03;
			14'd3352: ff_rdata <= 8'h30;
			14'd3353: ff_rdata <= 8'h70;
			14'd3354: ff_rdata <= 8'h19;
			14'd3355: ff_rdata <= 8'h20;
			14'd3356: ff_rdata <= 8'h42;
			14'd3357: ff_rdata <= 8'h62;
			14'd3358: ff_rdata <= 8'h26;
			14'd3359: ff_rdata <= 8'h24;
			14'd3360: ff_rdata <= 8'h62;
			14'd3361: ff_rdata <= 8'h71;
			14'd3362: ff_rdata <= 8'h25;
			14'd3363: ff_rdata <= 8'h20;
			14'd3364: ff_rdata <= 8'h64;
			14'd3365: ff_rdata <= 8'h43;
			14'd3366: ff_rdata <= 8'h12;
			14'd3367: ff_rdata <= 8'h26;
			14'd3368: ff_rdata <= 8'h21;
			14'd3369: ff_rdata <= 8'h03;
			14'd3370: ff_rdata <= 8'h0B;
			14'd3371: ff_rdata <= 8'h20;
			14'd3372: ff_rdata <= 8'h90;
			14'd3373: ff_rdata <= 8'hD4;
			14'd3374: ff_rdata <= 8'h02;
			14'd3375: ff_rdata <= 8'hF5;
			14'd3376: ff_rdata <= 8'h01;
			14'd3377: ff_rdata <= 8'h03;
			14'd3378: ff_rdata <= 8'h0A;
			14'd3379: ff_rdata <= 8'h20;
			14'd3380: ff_rdata <= 8'h90;
			14'd3381: ff_rdata <= 8'hA4;
			14'd3382: ff_rdata <= 8'h03;
			14'd3383: ff_rdata <= 8'hF5;
			14'd3384: ff_rdata <= 8'h43;
			14'd3385: ff_rdata <= 8'h53;
			14'd3386: ff_rdata <= 8'h0E;
			14'd3387: ff_rdata <= 8'h20;
			14'd3388: ff_rdata <= 8'hB5;
			14'd3389: ff_rdata <= 8'hE9;
			14'd3390: ff_rdata <= 8'h84;
			14'd3391: ff_rdata <= 8'h04;
			14'd3392: ff_rdata <= 8'h34;
			14'd3393: ff_rdata <= 8'h30;
			14'd3394: ff_rdata <= 8'h26;
			14'd3395: ff_rdata <= 8'h20;
			14'd3396: ff_rdata <= 8'h50;
			14'd3397: ff_rdata <= 8'h30;
			14'd3398: ff_rdata <= 8'h76;
			14'd3399: ff_rdata <= 8'h06;
			14'd3400: ff_rdata <= 8'h73;
			14'd3401: ff_rdata <= 8'h33;
			14'd3402: ff_rdata <= 8'h5A;
			14'd3403: ff_rdata <= 8'h20;
			14'd3404: ff_rdata <= 8'h99;
			14'd3405: ff_rdata <= 8'hF5;
			14'd3406: ff_rdata <= 8'h14;
			14'd3407: ff_rdata <= 8'h15;
			14'd3408: ff_rdata <= 8'h73;
			14'd3409: ff_rdata <= 8'h13;
			14'd3410: ff_rdata <= 8'h16;
			14'd3411: ff_rdata <= 8'h20;
			14'd3412: ff_rdata <= 8'hF9;
			14'd3413: ff_rdata <= 8'hF5;
			14'd3414: ff_rdata <= 8'h33;
			14'd3415: ff_rdata <= 8'h03;
			14'd3416: ff_rdata <= 8'h61;
			14'd3417: ff_rdata <= 8'h21;
			14'd3418: ff_rdata <= 8'h15;
			14'd3419: ff_rdata <= 8'h20;
			14'd3420: ff_rdata <= 8'h76;
			14'd3421: ff_rdata <= 8'h54;
			14'd3422: ff_rdata <= 8'h23;
			14'd3423: ff_rdata <= 8'h06;
			14'd3424: ff_rdata <= 8'h63;
			14'd3425: ff_rdata <= 8'h70;
			14'd3426: ff_rdata <= 8'h1B;
			14'd3427: ff_rdata <= 8'h20;
			14'd3428: ff_rdata <= 8'h75;
			14'd3429: ff_rdata <= 8'h4B;
			14'd3430: ff_rdata <= 8'h45;
			14'd3431: ff_rdata <= 8'h15;
			14'd3432: ff_rdata <= 8'h61;
			14'd3433: ff_rdata <= 8'hA1;
			14'd3434: ff_rdata <= 8'h0A;
			14'd3435: ff_rdata <= 8'h20;
			14'd3436: ff_rdata <= 8'h76;
			14'd3437: ff_rdata <= 8'h54;
			14'd3438: ff_rdata <= 8'h12;
			14'd3439: ff_rdata <= 8'h07;
			14'd3440: ff_rdata <= 8'h61;
			14'd3441: ff_rdata <= 8'h78;
			14'd3442: ff_rdata <= 8'h0D;
			14'd3443: ff_rdata <= 8'h20;
			14'd3444: ff_rdata <= 8'h85;
			14'd3445: ff_rdata <= 8'hF2;
			14'd3446: ff_rdata <= 8'h14;
			14'd3447: ff_rdata <= 8'h03;
			14'd3448: ff_rdata <= 8'h31;
			14'd3449: ff_rdata <= 8'h71;
			14'd3450: ff_rdata <= 8'h15;
			14'd3451: ff_rdata <= 8'h20;
			14'd3452: ff_rdata <= 8'hB6;
			14'd3453: ff_rdata <= 8'hF9;
			14'd3454: ff_rdata <= 8'h03;
			14'd3455: ff_rdata <= 8'h26;
			14'd3456: ff_rdata <= 8'h61;
			14'd3457: ff_rdata <= 8'h71;
			14'd3458: ff_rdata <= 8'h0D;
			14'd3459: ff_rdata <= 8'h20;
			14'd3460: ff_rdata <= 8'h75;
			14'd3461: ff_rdata <= 8'hF2;
			14'd3462: ff_rdata <= 8'h18;
			14'd3463: ff_rdata <= 8'h03;
			14'd3464: ff_rdata <= 8'h03;
			14'd3465: ff_rdata <= 8'h0C;
			14'd3466: ff_rdata <= 8'h14;
			14'd3467: ff_rdata <= 8'h20;
			14'd3468: ff_rdata <= 8'hA7;
			14'd3469: ff_rdata <= 8'hFC;
			14'd3470: ff_rdata <= 8'h13;
			14'd3471: ff_rdata <= 8'h15;
			14'd3472: ff_rdata <= 8'h13;
			14'd3473: ff_rdata <= 8'h32;
			14'd3474: ff_rdata <= 8'h80;
			14'd3475: ff_rdata <= 8'h20;
			14'd3476: ff_rdata <= 8'h20;
			14'd3477: ff_rdata <= 8'h85;
			14'd3478: ff_rdata <= 8'h03;
			14'd3479: ff_rdata <= 8'hAF;
			14'd3480: ff_rdata <= 8'hF1;
			14'd3481: ff_rdata <= 8'h31;
			14'd3482: ff_rdata <= 8'h17;
			14'd3483: ff_rdata <= 8'h20;
			14'd3484: ff_rdata <= 8'h23;
			14'd3485: ff_rdata <= 8'h40;
			14'd3486: ff_rdata <= 8'h14;
			14'd3487: ff_rdata <= 8'h09;
			14'd3488: ff_rdata <= 8'hF0;
			14'd3489: ff_rdata <= 8'h74;
			14'd3490: ff_rdata <= 8'h17;
			14'd3491: ff_rdata <= 8'h20;
			14'd3492: ff_rdata <= 8'h5A;
			14'd3493: ff_rdata <= 8'h43;
			14'd3494: ff_rdata <= 8'h06;
			14'd3495: ff_rdata <= 8'hFC;
			14'd3496: ff_rdata <= 8'h20;
			14'd3497: ff_rdata <= 8'h71;
			14'd3498: ff_rdata <= 8'h0D;
			14'd3499: ff_rdata <= 8'h20;
			14'd3500: ff_rdata <= 8'hC1;
			14'd3501: ff_rdata <= 8'hD5;
			14'd3502: ff_rdata <= 8'h56;
			14'd3503: ff_rdata <= 8'h06;
			14'd3504: ff_rdata <= 8'h30;
			14'd3505: ff_rdata <= 8'h32;
			14'd3506: ff_rdata <= 8'h06;
			14'd3507: ff_rdata <= 8'h20;
			14'd3508: ff_rdata <= 8'h40;
			14'd3509: ff_rdata <= 8'h40;
			14'd3510: ff_rdata <= 8'h04;
			14'd3511: ff_rdata <= 8'h74;
			14'd3512: ff_rdata <= 8'h30;
			14'd3513: ff_rdata <= 8'h32;
			14'd3514: ff_rdata <= 8'h03;
			14'd3515: ff_rdata <= 8'h20;
			14'd3516: ff_rdata <= 8'h40;
			14'd3517: ff_rdata <= 8'h40;
			14'd3518: ff_rdata <= 8'h04;
			14'd3519: ff_rdata <= 8'h74;
			14'd3520: ff_rdata <= 8'h01;
			14'd3521: ff_rdata <= 8'h08;
			14'd3522: ff_rdata <= 8'h0D;
			14'd3523: ff_rdata <= 8'h20;
			14'd3524: ff_rdata <= 8'h78;
			14'd3525: ff_rdata <= 8'hF8;
			14'd3526: ff_rdata <= 8'h7F;
			14'd3527: ff_rdata <= 8'hF9;
			14'd3528: ff_rdata <= 8'hC8;
			14'd3529: ff_rdata <= 8'hC0;
			14'd3530: ff_rdata <= 8'h0B;
			14'd3531: ff_rdata <= 8'h20;
			14'd3532: ff_rdata <= 8'h76;
			14'd3533: ff_rdata <= 8'hF7;
			14'd3534: ff_rdata <= 8'h11;
			14'd3535: ff_rdata <= 8'hF9;
			14'd3536: ff_rdata <= 8'h49;
			14'd3537: ff_rdata <= 8'h40;
			14'd3538: ff_rdata <= 8'h0B;
			14'd3539: ff_rdata <= 8'h20;
			14'd3540: ff_rdata <= 8'hB4;
			14'd3541: ff_rdata <= 8'hF9;
			14'd3542: ff_rdata <= 8'hFF;
			14'd3543: ff_rdata <= 8'h05;
			14'd3544: ff_rdata <= 8'hCD;
			14'd3545: ff_rdata <= 8'h42;
			14'd3546: ff_rdata <= 8'h0C;
			14'd3547: ff_rdata <= 8'h20;
			14'd3548: ff_rdata <= 8'hA2;
			14'd3549: ff_rdata <= 8'hF0;
			14'd3550: ff_rdata <= 8'h00;
			14'd3551: ff_rdata <= 8'h01;
			14'd3552: ff_rdata <= 8'h51;
			14'd3553: ff_rdata <= 8'h42;
			14'd3554: ff_rdata <= 8'h13;
			14'd3555: ff_rdata <= 8'h20;
			14'd3556: ff_rdata <= 8'h13;
			14'd3557: ff_rdata <= 8'h10;
			14'd3558: ff_rdata <= 8'h42;
			14'd3559: ff_rdata <= 8'h01;
			14'd3560: ff_rdata <= 8'h51;
			14'd3561: ff_rdata <= 8'h42;
			14'd3562: ff_rdata <= 8'h13;
			14'd3563: ff_rdata <= 8'h20;
			14'd3564: ff_rdata <= 8'h13;
			14'd3565: ff_rdata <= 8'h10;
			14'd3566: ff_rdata <= 8'h42;
			14'd3567: ff_rdata <= 8'h01;
			14'd3568: ff_rdata <= 8'h30;
			14'd3569: ff_rdata <= 8'h34;
			14'd3570: ff_rdata <= 8'h12;
			14'd3571: ff_rdata <= 8'h20;
			14'd3572: ff_rdata <= 8'h23;
			14'd3573: ff_rdata <= 8'h70;
			14'd3574: ff_rdata <= 8'h26;
			14'd3575: ff_rdata <= 8'h02;
			14'd3576: ff_rdata <= 8'h00;
			14'd3577: ff_rdata <= 8'h00;
			14'd3578: ff_rdata <= 8'hFF;
			14'd3579: ff_rdata <= 8'h20;
			14'd3580: ff_rdata <= 8'h00;
			14'd3581: ff_rdata <= 8'h00;
			14'd3582: ff_rdata <= 8'hFF;
			14'd3583: ff_rdata <= 8'hFF;
			14'd3584: ff_rdata <= 8'h21;
			14'd3585: ff_rdata <= 8'h00;
			14'd3586: ff_rdata <= 8'h00;
			14'd3587: ff_rdata <= 8'h00;
			14'd3588: ff_rdata <= 8'h00;
			14'd3589: ff_rdata <= 8'h00;
			14'd3590: ff_rdata <= 8'h00;
			14'd3591: ff_rdata <= 8'h00;
			14'd3592: ff_rdata <= 8'h00;
			14'd3593: ff_rdata <= 8'h00;
			14'd3594: ff_rdata <= 8'h00;
			14'd3595: ff_rdata <= 8'h00;
			14'd3596: ff_rdata <= 8'h00;
			14'd3597: ff_rdata <= 8'h00;
			14'd3598: ff_rdata <= 8'h00;
			14'd3599: ff_rdata <= 8'h00;
			14'd3600: ff_rdata <= 8'hB0;
			14'd3601: ff_rdata <= 8'h00;
			14'd3602: ff_rdata <= 8'h00;
			14'd3603: ff_rdata <= 8'h00;
			14'd3604: ff_rdata <= 8'h00;
			14'd3605: ff_rdata <= 8'h00;
			14'd3606: ff_rdata <= 8'h00;
			14'd3607: ff_rdata <= 8'h00;
			14'd3608: ff_rdata <= 8'h00;
			14'd3609: ff_rdata <= 8'h00;
			14'd3610: ff_rdata <= 8'h00;
			14'd3611: ff_rdata <= 8'h00;
			14'd3612: ff_rdata <= 8'h00;
			14'd3613: ff_rdata <= 8'h00;
			14'd3614: ff_rdata <= 8'h00;
			14'd3615: ff_rdata <= 8'h00;
			14'd3616: ff_rdata <= 8'h00;
			14'd3617: ff_rdata <= 8'h00;
			14'd3618: ff_rdata <= 8'h00;
			14'd3619: ff_rdata <= 8'h00;
			14'd3620: ff_rdata <= 8'h00;
			14'd3621: ff_rdata <= 8'h00;
			14'd3622: ff_rdata <= 8'h00;
			14'd3623: ff_rdata <= 8'h00;
			14'd3624: ff_rdata <= 8'h00;
			14'd3625: ff_rdata <= 8'hB3;
			14'd3626: ff_rdata <= 8'h00;
			14'd3627: ff_rdata <= 8'h00;
			14'd3628: ff_rdata <= 8'h00;
			14'd3629: ff_rdata <= 8'h00;
			14'd3630: ff_rdata <= 8'h00;
			14'd3631: ff_rdata <= 8'h00;
			14'd3632: ff_rdata <= 8'h00;
			14'd3633: ff_rdata <= 8'h00;
			14'd3634: ff_rdata <= 8'h00;
			14'd3635: ff_rdata <= 8'h00;
			14'd3636: ff_rdata <= 8'h00;
			14'd3637: ff_rdata <= 8'h00;
			14'd3638: ff_rdata <= 8'h00;
			14'd3639: ff_rdata <= 8'h00;
			14'd3640: ff_rdata <= 8'h00;
			14'd3641: ff_rdata <= 8'h00;
			14'd3642: ff_rdata <= 8'h00;
			14'd3643: ff_rdata <= 8'h00;
			14'd3644: ff_rdata <= 8'h00;
			14'd3645: ff_rdata <= 8'h00;
			14'd3646: ff_rdata <= 8'h00;
			14'd3647: ff_rdata <= 8'h00;
			14'd3648: ff_rdata <= 8'hFF;
			14'd3649: ff_rdata <= 8'hFF;
			14'd3650: ff_rdata <= 8'hB6;
			14'd3651: ff_rdata <= 8'hFF;
			14'd3652: ff_rdata <= 8'hFF;
			14'd3653: ff_rdata <= 8'hFF;
			14'd3654: ff_rdata <= 8'hFF;
			14'd3655: ff_rdata <= 8'hFF;
			14'd3656: ff_rdata <= 8'hFF;
			14'd3657: ff_rdata <= 8'hFF;
			14'd3658: ff_rdata <= 8'hFF;
			14'd3659: ff_rdata <= 8'hFF;
			14'd3660: ff_rdata <= 8'hFF;
			14'd3661: ff_rdata <= 8'hFF;
			14'd3662: ff_rdata <= 8'hFF;
			14'd3663: ff_rdata <= 8'hFF;
			14'd3664: ff_rdata <= 8'hFF;
			14'd3665: ff_rdata <= 8'hFF;
			14'd3666: ff_rdata <= 8'hFF;
			14'd3667: ff_rdata <= 8'hFF;
			14'd3668: ff_rdata <= 8'hFF;
			14'd3669: ff_rdata <= 8'hFF;
			14'd3670: ff_rdata <= 8'hFF;
			14'd3671: ff_rdata <= 8'hFF;
			14'd3672: ff_rdata <= 8'hFF;
			14'd3673: ff_rdata <= 8'hFF;
			14'd3674: ff_rdata <= 8'hFF;
			14'd3675: ff_rdata <= 8'hB9;
			14'd3676: ff_rdata <= 8'hFF;
			14'd3677: ff_rdata <= 8'hFF;
			14'd3678: ff_rdata <= 8'hFF;
			14'd3679: ff_rdata <= 8'hFF;
			14'd3680: ff_rdata <= 8'hFF;
			14'd3681: ff_rdata <= 8'hFF;
			14'd3682: ff_rdata <= 8'hFF;
			14'd3683: ff_rdata <= 8'hFF;
			14'd3684: ff_rdata <= 8'hFF;
			14'd3685: ff_rdata <= 8'hFF;
			14'd3686: ff_rdata <= 8'hFF;
			14'd3687: ff_rdata <= 8'hFF;
			14'd3688: ff_rdata <= 8'hFF;
			14'd3689: ff_rdata <= 8'hFF;
			14'd3690: ff_rdata <= 8'hFF;
			14'd3691: ff_rdata <= 8'hFF;
			14'd3692: ff_rdata <= 8'hFF;
			14'd3693: ff_rdata <= 8'hFF;
			14'd3694: ff_rdata <= 8'hFF;
			14'd3695: ff_rdata <= 8'hFF;
			14'd3696: ff_rdata <= 8'hFF;
			14'd3697: ff_rdata <= 8'hFF;
			14'd3698: ff_rdata <= 8'hFF;
			14'd3699: ff_rdata <= 8'hFF;
			14'd3700: ff_rdata <= 8'hBC;
			14'd3701: ff_rdata <= 8'hFF;
			14'd3702: ff_rdata <= 8'hFF;
			14'd3703: ff_rdata <= 8'hFF;
			14'd3704: ff_rdata <= 8'hFF;
			14'd3705: ff_rdata <= 8'hFF;
			14'd3706: ff_rdata <= 8'hFF;
			14'd3707: ff_rdata <= 8'hFF;
			14'd3708: ff_rdata <= 8'hFF;
			14'd3709: ff_rdata <= 8'hFF;
			14'd3710: ff_rdata <= 8'hFF;
			14'd3711: ff_rdata <= 8'h37;
			14'd3712: ff_rdata <= 8'h01;
			14'd3713: ff_rdata <= 8'h00;
			14'd3714: ff_rdata <= 8'h00;
			14'd3715: ff_rdata <= 8'h00;
			14'd3716: ff_rdata <= 8'h00;
			14'd3717: ff_rdata <= 8'h00;
			14'd3718: ff_rdata <= 8'h00;
			14'd3719: ff_rdata <= 8'h00;
			14'd3720: ff_rdata <= 8'h00;
			14'd3721: ff_rdata <= 8'h00;
			14'd3722: ff_rdata <= 8'h00;
			14'd3723: ff_rdata <= 8'h00;
			14'd3724: ff_rdata <= 8'h00;
			14'd3725: ff_rdata <= 8'hBF;
			14'd3726: ff_rdata <= 8'h00;
			14'd3727: ff_rdata <= 8'h00;
			14'd3728: ff_rdata <= 8'h00;
			14'd3729: ff_rdata <= 8'h00;
			14'd3730: ff_rdata <= 8'h00;
			14'd3731: ff_rdata <= 8'h00;
			14'd3732: ff_rdata <= 8'h00;
			14'd3733: ff_rdata <= 8'h00;
			14'd3734: ff_rdata <= 8'h00;
			14'd3735: ff_rdata <= 8'h00;
			14'd3736: ff_rdata <= 8'h00;
			14'd3737: ff_rdata <= 8'h00;
			14'd3738: ff_rdata <= 8'h00;
			14'd3739: ff_rdata <= 8'h00;
			14'd3740: ff_rdata <= 8'h00;
			14'd3741: ff_rdata <= 8'h00;
			14'd3742: ff_rdata <= 8'h00;
			14'd3743: ff_rdata <= 8'h00;
			14'd3744: ff_rdata <= 8'h00;
			14'd3745: ff_rdata <= 8'h00;
			14'd3746: ff_rdata <= 8'h00;
			14'd3747: ff_rdata <= 8'h00;
			14'd3748: ff_rdata <= 8'h00;
			14'd3749: ff_rdata <= 8'h00;
			14'd3750: ff_rdata <= 8'hC2;
			14'd3751: ff_rdata <= 8'h00;
			14'd3752: ff_rdata <= 8'h00;
			14'd3753: ff_rdata <= 8'h00;
			14'd3754: ff_rdata <= 8'h00;
			14'd3755: ff_rdata <= 8'h00;
			14'd3756: ff_rdata <= 8'h00;
			14'd3757: ff_rdata <= 8'h00;
			14'd3758: ff_rdata <= 8'h00;
			14'd3759: ff_rdata <= 8'h00;
			14'd3760: ff_rdata <= 8'h00;
			14'd3761: ff_rdata <= 8'h00;
			14'd3762: ff_rdata <= 8'h00;
			14'd3763: ff_rdata <= 8'h00;
			14'd3764: ff_rdata <= 8'h00;
			14'd3765: ff_rdata <= 8'h00;
			14'd3766: ff_rdata <= 8'h00;
			14'd3767: ff_rdata <= 8'h00;
			14'd3768: ff_rdata <= 8'h00;
			14'd3769: ff_rdata <= 8'h00;
			14'd3770: ff_rdata <= 8'h00;
			14'd3771: ff_rdata <= 8'h00;
			14'd3772: ff_rdata <= 8'h00;
			14'd3773: ff_rdata <= 8'h00;
			14'd3774: ff_rdata <= 8'h00;
			14'd3775: ff_rdata <= 8'hC5;
			14'd3776: ff_rdata <= 8'hFF;
			14'd3777: ff_rdata <= 8'hFF;
			14'd3778: ff_rdata <= 8'hFF;
			14'd3779: ff_rdata <= 8'hFF;
			14'd3780: ff_rdata <= 8'hFF;
			14'd3781: ff_rdata <= 8'hFF;
			14'd3782: ff_rdata <= 8'hFF;
			14'd3783: ff_rdata <= 8'hFF;
			14'd3784: ff_rdata <= 8'hFF;
			14'd3785: ff_rdata <= 8'hFF;
			14'd3786: ff_rdata <= 8'hFF;
			14'd3787: ff_rdata <= 8'hFF;
			14'd3788: ff_rdata <= 8'hFF;
			14'd3789: ff_rdata <= 8'hFF;
			14'd3790: ff_rdata <= 8'hFF;
			14'd3791: ff_rdata <= 8'hFF;
			14'd3792: ff_rdata <= 8'hFF;
			14'd3793: ff_rdata <= 8'hFF;
			14'd3794: ff_rdata <= 8'hFF;
			14'd3795: ff_rdata <= 8'hFF;
			14'd3796: ff_rdata <= 8'hFF;
			14'd3797: ff_rdata <= 8'hFF;
			14'd3798: ff_rdata <= 8'hFF;
			14'd3799: ff_rdata <= 8'hFF;
			14'd3800: ff_rdata <= 8'hC8;
			14'd3801: ff_rdata <= 8'hFF;
			14'd3802: ff_rdata <= 8'hFF;
			14'd3803: ff_rdata <= 8'hFF;
			14'd3804: ff_rdata <= 8'hFF;
			14'd3805: ff_rdata <= 8'hFF;
			14'd3806: ff_rdata <= 8'hFF;
			14'd3807: ff_rdata <= 8'hFF;
			14'd3808: ff_rdata <= 8'hFF;
			14'd3809: ff_rdata <= 8'hFF;
			14'd3810: ff_rdata <= 8'hFF;
			14'd3811: ff_rdata <= 8'hFF;
			14'd3812: ff_rdata <= 8'hFF;
			14'd3813: ff_rdata <= 8'hFF;
			14'd3814: ff_rdata <= 8'hFF;
			14'd3815: ff_rdata <= 8'hFF;
			14'd3816: ff_rdata <= 8'hFF;
			14'd3817: ff_rdata <= 8'hFF;
			14'd3818: ff_rdata <= 8'hFF;
			14'd3819: ff_rdata <= 8'hFF;
			14'd3820: ff_rdata <= 8'hFF;
			14'd3821: ff_rdata <= 8'hFF;
			14'd3822: ff_rdata <= 8'hFF;
			14'd3823: ff_rdata <= 8'hFF;
			14'd3824: ff_rdata <= 8'hFF;
			14'd3825: ff_rdata <= 8'hCB;
			14'd3826: ff_rdata <= 8'hFF;
			14'd3827: ff_rdata <= 8'hFF;
			14'd3828: ff_rdata <= 8'hFF;
			14'd3829: ff_rdata <= 8'hFF;
			14'd3830: ff_rdata <= 8'hFF;
			14'd3831: ff_rdata <= 8'hFF;
			14'd3832: ff_rdata <= 8'hFF;
			14'd3833: ff_rdata <= 8'hFF;
			14'd3834: ff_rdata <= 8'hFF;
			14'd3835: ff_rdata <= 8'hFF;
			14'd3836: ff_rdata <= 8'hFF;
			14'd3837: ff_rdata <= 8'hFF;
			14'd3838: ff_rdata <= 8'hFF;
			14'd3839: ff_rdata <= 8'hFF;
			14'd3840: ff_rdata <= 8'hFF;
			14'd3841: ff_rdata <= 8'hFF;
			14'd3842: ff_rdata <= 8'hFF;
			14'd3843: ff_rdata <= 8'hFF;
			14'd3844: ff_rdata <= 8'hFF;
			14'd3845: ff_rdata <= 8'hFF;
			14'd3846: ff_rdata <= 8'hFF;
			14'd3847: ff_rdata <= 8'hFF;
			14'd3848: ff_rdata <= 8'hFF;
			14'd3849: ff_rdata <= 8'hFF;
			14'd3850: ff_rdata <= 8'hCE;
			14'd3851: ff_rdata <= 8'hFF;
			14'd3852: ff_rdata <= 8'hFF;
			14'd3853: ff_rdata <= 8'hFF;
			14'd3854: ff_rdata <= 8'hFF;
			14'd3855: ff_rdata <= 8'hFF;
			14'd3856: ff_rdata <= 8'hFF;
			14'd3857: ff_rdata <= 8'hFF;
			14'd3858: ff_rdata <= 8'hFF;
			14'd3859: ff_rdata <= 8'hFF;
			14'd3860: ff_rdata <= 8'hFF;
			14'd3861: ff_rdata <= 8'hFF;
			14'd3862: ff_rdata <= 8'hFF;
			14'd3863: ff_rdata <= 8'hFF;
			14'd3864: ff_rdata <= 8'hFF;
			14'd3865: ff_rdata <= 8'hFF;
			14'd3866: ff_rdata <= 8'hFF;
			14'd3867: ff_rdata <= 8'hFF;
			14'd3868: ff_rdata <= 8'hFF;
			14'd3869: ff_rdata <= 8'hFF;
			14'd3870: ff_rdata <= 8'hFF;
			14'd3871: ff_rdata <= 8'hFF;
			14'd3872: ff_rdata <= 8'hFF;
			14'd3873: ff_rdata <= 8'hFF;
			14'd3874: ff_rdata <= 8'hFF;
			14'd3875: ff_rdata <= 8'hD1;
			14'd3876: ff_rdata <= 8'hFF;
			14'd3877: ff_rdata <= 8'hFF;
			14'd3878: ff_rdata <= 8'hFF;
			14'd3879: ff_rdata <= 8'hFF;
			14'd3880: ff_rdata <= 8'hFF;
			14'd3881: ff_rdata <= 8'hFF;
			14'd3882: ff_rdata <= 8'hFF;
			14'd3883: ff_rdata <= 8'hFF;
			14'd3884: ff_rdata <= 8'hFF;
			14'd3885: ff_rdata <= 8'hFF;
			14'd3886: ff_rdata <= 8'hFF;
			14'd3887: ff_rdata <= 8'hFF;
			14'd3888: ff_rdata <= 8'hFF;
			14'd3889: ff_rdata <= 8'hFF;
			14'd3890: ff_rdata <= 8'hFF;
			14'd3891: ff_rdata <= 8'hFF;
			14'd3892: ff_rdata <= 8'hFF;
			14'd3893: ff_rdata <= 8'hFF;
			14'd3894: ff_rdata <= 8'hFF;
			14'd3895: ff_rdata <= 8'hFF;
			14'd3896: ff_rdata <= 8'hFF;
			14'd3897: ff_rdata <= 8'hFF;
			14'd3898: ff_rdata <= 8'hFF;
			14'd3899: ff_rdata <= 8'hFF;
			14'd3900: ff_rdata <= 8'hD4;
			14'd3901: ff_rdata <= 8'hFF;
			14'd3902: ff_rdata <= 8'hFF;
			14'd3903: ff_rdata <= 8'hFF;
			14'd3904: ff_rdata <= 8'h00;
			14'd3905: ff_rdata <= 8'h00;
			14'd3906: ff_rdata <= 8'h00;
			14'd3907: ff_rdata <= 8'h00;
			14'd3908: ff_rdata <= 8'h00;
			14'd3909: ff_rdata <= 8'h00;
			14'd3910: ff_rdata <= 8'h00;
			14'd3911: ff_rdata <= 8'h00;
			14'd3912: ff_rdata <= 8'h00;
			14'd3913: ff_rdata <= 8'h00;
			14'd3914: ff_rdata <= 8'h00;
			14'd3915: ff_rdata <= 8'h00;
			14'd3916: ff_rdata <= 8'h00;
			14'd3917: ff_rdata <= 8'h00;
			14'd3918: ff_rdata <= 8'h00;
			14'd3919: ff_rdata <= 8'h00;
			14'd3920: ff_rdata <= 8'h00;
			14'd3921: ff_rdata <= 8'h00;
			14'd3922: ff_rdata <= 8'h00;
			14'd3923: ff_rdata <= 8'h00;
			14'd3924: ff_rdata <= 8'h00;
			14'd3925: ff_rdata <= 8'hD7;
			14'd3926: ff_rdata <= 8'h00;
			14'd3927: ff_rdata <= 8'h00;
			14'd3928: ff_rdata <= 8'h00;
			14'd3929: ff_rdata <= 8'h00;
			14'd3930: ff_rdata <= 8'h00;
			14'd3931: ff_rdata <= 8'h00;
			14'd3932: ff_rdata <= 8'h00;
			14'd3933: ff_rdata <= 8'h00;
			14'd3934: ff_rdata <= 8'h00;
			14'd3935: ff_rdata <= 8'h00;
			14'd3936: ff_rdata <= 8'h00;
			14'd3937: ff_rdata <= 8'h00;
			14'd3938: ff_rdata <= 8'h00;
			14'd3939: ff_rdata <= 8'h00;
			14'd3940: ff_rdata <= 8'h00;
			14'd3941: ff_rdata <= 8'h00;
			14'd3942: ff_rdata <= 8'h00;
			14'd3943: ff_rdata <= 8'h00;
			14'd3944: ff_rdata <= 8'h00;
			14'd3945: ff_rdata <= 8'h00;
			14'd3946: ff_rdata <= 8'h00;
			14'd3947: ff_rdata <= 8'h00;
			14'd3948: ff_rdata <= 8'h00;
			14'd3949: ff_rdata <= 8'h00;
			14'd3950: ff_rdata <= 8'hDA;
			14'd3951: ff_rdata <= 8'h00;
			14'd3952: ff_rdata <= 8'h00;
			14'd3953: ff_rdata <= 8'h00;
			14'd3954: ff_rdata <= 8'h00;
			14'd3955: ff_rdata <= 8'h00;
			14'd3956: ff_rdata <= 8'h00;
			14'd3957: ff_rdata <= 8'h00;
			14'd3958: ff_rdata <= 8'h00;
			14'd3959: ff_rdata <= 8'h00;
			14'd3960: ff_rdata <= 8'h00;
			14'd3961: ff_rdata <= 8'h00;
			14'd3962: ff_rdata <= 8'h00;
			14'd3963: ff_rdata <= 8'h00;
			14'd3964: ff_rdata <= 8'h00;
			14'd3965: ff_rdata <= 8'h00;
			14'd3966: ff_rdata <= 8'h00;
			14'd3967: ff_rdata <= 8'hC9;
			14'd3968: ff_rdata <= 8'hDF;
			14'd3969: ff_rdata <= 8'hFF;
			14'd3970: ff_rdata <= 8'hFF;
			14'd3971: ff_rdata <= 8'hFF;
			14'd3972: ff_rdata <= 8'hFF;
			14'd3973: ff_rdata <= 8'hFF;
			14'd3974: ff_rdata <= 8'hFF;
			14'd3975: ff_rdata <= 8'hDD;
			14'd3976: ff_rdata <= 8'hFF;
			14'd3977: ff_rdata <= 8'hFF;
			14'd3978: ff_rdata <= 8'hFF;
			14'd3979: ff_rdata <= 8'hFF;
			14'd3980: ff_rdata <= 8'hFF;
			14'd3981: ff_rdata <= 8'hFF;
			14'd3982: ff_rdata <= 8'hFF;
			14'd3983: ff_rdata <= 8'hFF;
			14'd3984: ff_rdata <= 8'hFF;
			14'd3985: ff_rdata <= 8'hFF;
			14'd3986: ff_rdata <= 8'hFF;
			14'd3987: ff_rdata <= 8'hFF;
			14'd3988: ff_rdata <= 8'hFF;
			14'd3989: ff_rdata <= 8'hFF;
			14'd3990: ff_rdata <= 8'hFF;
			14'd3991: ff_rdata <= 8'hFF;
			14'd3992: ff_rdata <= 8'hFF;
			14'd3993: ff_rdata <= 8'hFF;
			14'd3994: ff_rdata <= 8'hFF;
			14'd3995: ff_rdata <= 8'hFF;
			14'd3996: ff_rdata <= 8'hFF;
			14'd3997: ff_rdata <= 8'hFF;
			14'd3998: ff_rdata <= 8'hFF;
			14'd3999: ff_rdata <= 8'hFF;
			14'd4000: ff_rdata <= 8'hE0;
			14'd4001: ff_rdata <= 8'hFF;
			14'd4002: ff_rdata <= 8'hFF;
			14'd4003: ff_rdata <= 8'hFF;
			14'd4004: ff_rdata <= 8'hFF;
			14'd4005: ff_rdata <= 8'hFF;
			14'd4006: ff_rdata <= 8'hFF;
			14'd4007: ff_rdata <= 8'hFF;
			14'd4008: ff_rdata <= 8'hFF;
			14'd4009: ff_rdata <= 8'hFF;
			14'd4010: ff_rdata <= 8'hFF;
			14'd4011: ff_rdata <= 8'hFF;
			14'd4012: ff_rdata <= 8'hFF;
			14'd4013: ff_rdata <= 8'hFF;
			14'd4014: ff_rdata <= 8'hFF;
			14'd4015: ff_rdata <= 8'hFF;
			14'd4016: ff_rdata <= 8'hFF;
			14'd4017: ff_rdata <= 8'hFF;
			14'd4018: ff_rdata <= 8'hFF;
			14'd4019: ff_rdata <= 8'hFF;
			14'd4020: ff_rdata <= 8'hFF;
			14'd4021: ff_rdata <= 8'hFF;
			14'd4022: ff_rdata <= 8'hFF;
			14'd4023: ff_rdata <= 8'hFF;
			14'd4024: ff_rdata <= 8'hFF;
			14'd4025: ff_rdata <= 8'hE3;
			14'd4026: ff_rdata <= 8'hFF;
			14'd4027: ff_rdata <= 8'hFF;
			14'd4028: ff_rdata <= 8'hFF;
			14'd4029: ff_rdata <= 8'hFF;
			14'd4030: ff_rdata <= 8'hFF;
			14'd4031: ff_rdata <= 8'hFF;
			14'd4032: ff_rdata <= 8'h00;
			14'd4033: ff_rdata <= 8'h00;
			14'd4034: ff_rdata <= 8'h00;
			14'd4035: ff_rdata <= 8'h00;
			14'd4036: ff_rdata <= 8'h00;
			14'd4037: ff_rdata <= 8'h00;
			14'd4038: ff_rdata <= 8'h00;
			14'd4039: ff_rdata <= 8'h00;
			14'd4040: ff_rdata <= 8'h00;
			14'd4041: ff_rdata <= 8'h00;
			14'd4042: ff_rdata <= 8'h00;
			14'd4043: ff_rdata <= 8'h00;
			14'd4044: ff_rdata <= 8'h00;
			14'd4045: ff_rdata <= 8'h00;
			14'd4046: ff_rdata <= 8'h00;
			14'd4047: ff_rdata <= 8'h00;
			14'd4048: ff_rdata <= 8'h00;
			14'd4049: ff_rdata <= 8'h00;
			14'd4050: ff_rdata <= 8'hE6;
			14'd4051: ff_rdata <= 8'h00;
			14'd4052: ff_rdata <= 8'h00;
			14'd4053: ff_rdata <= 8'h00;
			14'd4054: ff_rdata <= 8'h00;
			14'd4055: ff_rdata <= 8'h00;
			14'd4056: ff_rdata <= 8'h00;
			14'd4057: ff_rdata <= 8'h00;
			14'd4058: ff_rdata <= 8'h00;
			14'd4059: ff_rdata <= 8'h00;
			14'd4060: ff_rdata <= 8'h00;
			14'd4061: ff_rdata <= 8'h00;
			14'd4062: ff_rdata <= 8'h00;
			14'd4063: ff_rdata <= 8'h00;
			14'd4064: ff_rdata <= 8'h00;
			14'd4065: ff_rdata <= 8'h00;
			14'd4066: ff_rdata <= 8'h00;
			14'd4067: ff_rdata <= 8'h00;
			14'd4068: ff_rdata <= 8'h00;
			14'd4069: ff_rdata <= 8'h00;
			14'd4070: ff_rdata <= 8'h00;
			14'd4071: ff_rdata <= 8'h00;
			14'd4072: ff_rdata <= 8'h00;
			14'd4073: ff_rdata <= 8'h00;
			14'd4074: ff_rdata <= 8'h00;
			14'd4075: ff_rdata <= 8'hE9;
			14'd4076: ff_rdata <= 8'h00;
			14'd4077: ff_rdata <= 8'h00;
			14'd4078: ff_rdata <= 8'h00;
			14'd4079: ff_rdata <= 8'h00;
			14'd4080: ff_rdata <= 8'h00;
			14'd4081: ff_rdata <= 8'h00;
			14'd4082: ff_rdata <= 8'h00;
			14'd4083: ff_rdata <= 8'h00;
			14'd4084: ff_rdata <= 8'h00;
			14'd4085: ff_rdata <= 8'h00;
			14'd4086: ff_rdata <= 8'h00;
			14'd4087: ff_rdata <= 8'h00;
			14'd4088: ff_rdata <= 8'h00;
			14'd4089: ff_rdata <= 8'h00;
			14'd4090: ff_rdata <= 8'h00;
			14'd4091: ff_rdata <= 8'h00;
			14'd4092: ff_rdata <= 8'h00;
			14'd4093: ff_rdata <= 8'h00;
			14'd4094: ff_rdata <= 8'h00;
			14'd4095: ff_rdata <= 8'h00;
			14'd4096: ff_rdata <= 8'hC3;
			14'd4097: ff_rdata <= 8'hEB;
			14'd4098: ff_rdata <= 8'h50;
			14'd4099: ff_rdata <= 8'hC3;
			14'd4100: ff_rdata <= 8'h5B;
			14'd4101: ff_rdata <= 8'h60;
			14'd4102: ff_rdata <= 8'hC3;
			14'd4103: ff_rdata <= 8'h78;
			14'd4104: ff_rdata <= 8'h50;
			14'd4105: ff_rdata <= 8'h21;
			14'd4106: ff_rdata <= 8'h75;
			14'd4107: ff_rdata <= 8'hF9;
			14'd4108: ff_rdata <= 8'h11;
			14'd4109: ff_rdata <= 8'h76;
			14'd4110: ff_rdata <= 8'hF9;
			14'd4111: ff_rdata <= 8'h01;
			14'd4112: ff_rdata <= 8'h46;
			14'd4113: ff_rdata <= 8'h01;
			14'd4114: ff_rdata <= 8'h36;
			14'd4115: ff_rdata <= 8'h00;
			14'd4116: ff_rdata <= 8'hED;
			14'd4117: ff_rdata <= 8'hB0;
			14'd4118: ff_rdata <= 8'h06;
			14'd4119: ff_rdata <= 8'h04;
			14'd4120: ff_rdata <= 8'hC5;
			14'd4121: ff_rdata <= 8'h3E;
			14'd4122: ff_rdata <= 8'h04;
			14'd4123: ff_rdata <= 8'h90;
			14'd4124: ff_rdata <= 8'h4F;
			14'd4125: ff_rdata <= 8'h21;
			14'd4126: ff_rdata <= 8'hC1;
			14'd4127: ff_rdata <= 8'hFC;
			14'd4128: ff_rdata <= 8'hCD;
			14'd4129: ff_rdata <= 8'h86;
			14'd4130: ff_rdata <= 8'h54;
			14'd4131: ff_rdata <= 8'h7E;
			14'd4132: ff_rdata <= 8'h87;
			14'd4133: ff_rdata <= 8'h30;
			14'd4134: ff_rdata <= 8'h1C;
			14'd4135: ff_rdata <= 8'h06;
			14'd4136: ff_rdata <= 8'h04;
			14'd4137: ff_rdata <= 8'hC5;
			14'd4138: ff_rdata <= 8'h3E;
			14'd4139: ff_rdata <= 8'h24;
			14'd4140: ff_rdata <= 8'h90;
			14'd4141: ff_rdata <= 8'h07;
			14'd4142: ff_rdata <= 8'h07;
			14'd4143: ff_rdata <= 8'hB1;
			14'd4144: ff_rdata <= 8'hCD;
			14'd4145: ff_rdata <= 8'h54;
			14'd4146: ff_rdata <= 8'h50;
			14'd4147: ff_rdata <= 8'hC1;
			14'd4148: ff_rdata <= 8'h28;
			14'd4149: ff_rdata <= 8'h13;
			14'd4150: ff_rdata <= 8'h10;
			14'd4151: ff_rdata <= 8'hF1;
			14'd4152: ff_rdata <= 8'hC1;
			14'd4153: ff_rdata <= 8'h10;
			14'd4154: ff_rdata <= 8'hDD;
			14'd4155: ff_rdata <= 8'h21;
			14'd4156: ff_rdata <= 8'hF6;
			14'd4157: ff_rdata <= 8'h7F;
			14'd4158: ff_rdata <= 8'hCB;
			14'd4159: ff_rdata <= 8'hC6;
			14'd4160: ff_rdata <= 8'hC3;
			14'd4161: ff_rdata <= 8'h61;
			14'd4162: ff_rdata <= 8'h6D;
			14'd4163: ff_rdata <= 8'h79;
			14'd4164: ff_rdata <= 8'hCD;
			14'd4165: ff_rdata <= 8'h54;
			14'd4166: ff_rdata <= 8'h50;
			14'd4167: ff_rdata <= 8'h20;
			14'd4168: ff_rdata <= 8'hEF;
			14'd4169: ff_rdata <= 8'hC1;
			14'd4170: ff_rdata <= 8'h18;
			14'd4171: ff_rdata <= 8'hF4;
			14'd4172: ff_rdata <= 8'h41;
			14'd4173: ff_rdata <= 8'h50;
			14'd4174: ff_rdata <= 8'h52;
			14'd4175: ff_rdata <= 8'h4C;
			14'd4176: ff_rdata <= 8'h4F;
			14'd4177: ff_rdata <= 8'h50;
			14'd4178: ff_rdata <= 8'h4C;
			14'd4179: ff_rdata <= 8'h4C;
			14'd4180: ff_rdata <= 8'hC5;
			14'd4181: ff_rdata <= 8'h21;
			14'd4182: ff_rdata <= 8'h18;
			14'd4183: ff_rdata <= 8'h40;
			14'd4184: ff_rdata <= 8'h11;
			14'd4185: ff_rdata <= 8'h4C;
			14'd4186: ff_rdata <= 8'h50;
			14'd4187: ff_rdata <= 8'h06;
			14'd4188: ff_rdata <= 8'h08;
			14'd4189: ff_rdata <= 8'hF5;
			14'd4190: ff_rdata <= 8'hC5;
			14'd4191: ff_rdata <= 8'hD5;
			14'd4192: ff_rdata <= 8'hCD;
			14'd4193: ff_rdata <= 8'h0C;
			14'd4194: ff_rdata <= 8'h00;
			14'd4195: ff_rdata <= 8'hFB;
			14'd4196: ff_rdata <= 8'hD1;
			14'd4197: ff_rdata <= 8'hC1;
			14'd4198: ff_rdata <= 8'h4F;
			14'd4199: ff_rdata <= 8'h1A;
			14'd4200: ff_rdata <= 8'hB9;
			14'd4201: ff_rdata <= 8'h20;
			14'd4202: ff_rdata <= 8'h08;
			14'd4203: ff_rdata <= 8'hF1;
			14'd4204: ff_rdata <= 8'h13;
			14'd4205: ff_rdata <= 8'h23;
			14'd4206: ff_rdata <= 8'h10;
			14'd4207: ff_rdata <= 8'hED;
			14'd4208: ff_rdata <= 8'hC1;
			14'd4209: ff_rdata <= 8'hAF;
			14'd4210: ff_rdata <= 8'hC9;
			14'd4211: ff_rdata <= 8'hF1;
			14'd4212: ff_rdata <= 8'hC1;
			14'd4213: ff_rdata <= 8'hAF;
			14'd4214: ff_rdata <= 8'h3C;
			14'd4215: ff_rdata <= 8'hC9;
			14'd4216: ff_rdata <= 8'hCD;
			14'd4217: ff_rdata <= 8'hC6;
			14'd4218: ff_rdata <= 8'h50;
			14'd4219: ff_rdata <= 8'hC8;
			14'd4220: ff_rdata <= 8'hC3;
			14'd4221: ff_rdata <= 8'h8D;
			14'd4222: ff_rdata <= 8'h65;
			14'd4223: ff_rdata <= 8'hF3;
			14'd4224: ff_rdata <= 8'hCD;
			14'd4225: ff_rdata <= 8'hC6;
			14'd4226: ff_rdata <= 8'h50;
			14'd4227: ff_rdata <= 8'hC0;
			14'd4228: ff_rdata <= 8'hCD;
			14'd4229: ff_rdata <= 8'hBE;
			14'd4230: ff_rdata <= 8'h50;
			14'd4231: ff_rdata <= 8'h21;
			14'd4232: ff_rdata <= 8'h9F;
			14'd4233: ff_rdata <= 8'hFD;
			14'd4234: ff_rdata <= 8'h11;
			14'd4235: ff_rdata <= 8'hBB;
			14'd4236: ff_rdata <= 8'hF9;
			14'd4237: ff_rdata <= 8'hE5;
			14'd4238: ff_rdata <= 8'hCD;
			14'd4239: ff_rdata <= 8'hAE;
			14'd4240: ff_rdata <= 8'h50;
			14'd4241: ff_rdata <= 8'h21;
			14'd4242: ff_rdata <= 8'hB9;
			14'd4243: ff_rdata <= 8'h50;
			14'd4244: ff_rdata <= 8'hD1;
			14'd4245: ff_rdata <= 8'hCD;
			14'd4246: ff_rdata <= 8'hAE;
			14'd4247: ff_rdata <= 8'h50;
			14'd4248: ff_rdata <= 8'hCD;
			14'd4249: ff_rdata <= 8'h4C;
			14'd4250: ff_rdata <= 8'h55;
			14'd4251: ff_rdata <= 8'h32;
			14'd4252: ff_rdata <= 8'h7C;
			14'd4253: ff_rdata <= 8'hF9;
			14'd4254: ff_rdata <= 8'h32;
			14'd4255: ff_rdata <= 8'hA0;
			14'd4256: ff_rdata <= 8'hFD;
			14'd4257: ff_rdata <= 8'h21;
			14'd4258: ff_rdata <= 8'hB4;
			14'd4259: ff_rdata <= 8'h50;
			14'd4260: ff_rdata <= 8'h11;
			14'd4261: ff_rdata <= 8'hC5;
			14'd4262: ff_rdata <= 8'hFF;
			14'd4263: ff_rdata <= 8'hCD;
			14'd4264: ff_rdata <= 8'hAE;
			14'd4265: ff_rdata <= 8'h50;
			14'd4266: ff_rdata <= 8'h32;
			14'd4267: ff_rdata <= 8'hC6;
			14'd4268: ff_rdata <= 8'hFF;
			14'd4269: ff_rdata <= 8'hC9;
			14'd4270: ff_rdata <= 8'h01;
			14'd4271: ff_rdata <= 8'h05;
			14'd4272: ff_rdata <= 8'h00;
			14'd4273: ff_rdata <= 8'hED;
			14'd4274: ff_rdata <= 8'hB0;
			14'd4275: ff_rdata <= 8'hC9;
			14'd4276: ff_rdata <= 8'hF7;
			14'd4277: ff_rdata <= 8'h00;
			14'd4278: ff_rdata <= 8'hA1;
			14'd4279: ff_rdata <= 8'h57;
			14'd4280: ff_rdata <= 8'hC9;
			14'd4281: ff_rdata <= 8'hF7;
			14'd4282: ff_rdata <= 8'h00;
			14'd4283: ff_rdata <= 8'hED;
			14'd4284: ff_rdata <= 8'h7F;
			14'd4285: ff_rdata <= 8'hC9;
			14'd4286: ff_rdata <= 8'hE5;
			14'd4287: ff_rdata <= 8'hCD;
			14'd4288: ff_rdata <= 8'hCE;
			14'd4289: ff_rdata <= 8'h50;
			14'd4290: ff_rdata <= 8'hCB;
			14'd4291: ff_rdata <= 8'hC6;
			14'd4292: ff_rdata <= 8'hE1;
			14'd4293: ff_rdata <= 8'hC9;
			14'd4294: ff_rdata <= 8'hE5;
			14'd4295: ff_rdata <= 8'hCD;
			14'd4296: ff_rdata <= 8'hCE;
			14'd4297: ff_rdata <= 8'h50;
			14'd4298: ff_rdata <= 8'hCB;
			14'd4299: ff_rdata <= 8'h46;
			14'd4300: ff_rdata <= 8'hE1;
			14'd4301: ff_rdata <= 8'hC9;
			14'd4302: ff_rdata <= 8'hF5;
			14'd4303: ff_rdata <= 8'hD5;
			14'd4304: ff_rdata <= 8'hCD;
			14'd4305: ff_rdata <= 8'h4C;
			14'd4306: ff_rdata <= 8'h55;
			14'd4307: ff_rdata <= 8'hE6;
			14'd4308: ff_rdata <= 8'h0F;
			14'd4309: ff_rdata <= 8'h6F;
			14'd4310: ff_rdata <= 8'h07;
			14'd4311: ff_rdata <= 8'h07;
			14'd4312: ff_rdata <= 8'h07;
			14'd4313: ff_rdata <= 8'h07;
			14'd4314: ff_rdata <= 8'hE6;
			14'd4315: ff_rdata <= 8'h30;
			14'd4316: ff_rdata <= 8'hB5;
			14'd4317: ff_rdata <= 8'hE6;
			14'd4318: ff_rdata <= 8'h3C;
			14'd4319: ff_rdata <= 8'h3C;
			14'd4320: ff_rdata <= 8'h87;
			14'd4321: ff_rdata <= 8'h5F;
			14'd4322: ff_rdata <= 8'h16;
			14'd4323: ff_rdata <= 8'h00;
			14'd4324: ff_rdata <= 8'h21;
			14'd4325: ff_rdata <= 8'h09;
			14'd4326: ff_rdata <= 8'hFD;
			14'd4327: ff_rdata <= 8'h19;
			14'd4328: ff_rdata <= 8'hD1;
			14'd4329: ff_rdata <= 8'hF1;
			14'd4330: ff_rdata <= 8'hC9;
			14'd4331: ff_rdata <= 8'hFB;
			14'd4332: ff_rdata <= 8'hE5;
			14'd4333: ff_rdata <= 8'h21;
			14'd4334: ff_rdata <= 8'h89;
			14'd4335: ff_rdata <= 8'hFD;
			14'd4336: ff_rdata <= 8'hCD;
			14'd4337: ff_rdata <= 8'h5A;
			14'd4338: ff_rdata <= 8'h52;
			14'd4339: ff_rdata <= 8'hE1;
			14'd4340: ff_rdata <= 8'hD8;
			14'd4341: ff_rdata <= 8'hE5;
			14'd4342: ff_rdata <= 8'h21;
			14'd4343: ff_rdata <= 8'hEC;
			14'd4344: ff_rdata <= 8'h52;
			14'd4345: ff_rdata <= 8'hB7;
			14'd4346: ff_rdata <= 8'hED;
			14'd4347: ff_rdata <= 8'h52;
			14'd4348: ff_rdata <= 8'hE1;
			14'd4349: ff_rdata <= 8'h28;
			14'd4350: ff_rdata <= 8'h05;
			14'd4351: ff_rdata <= 8'hCD;
			14'd4352: ff_rdata <= 8'hC6;
			14'd4353: ff_rdata <= 8'h50;
			14'd4354: ff_rdata <= 8'h37;
			14'd4355: ff_rdata <= 8'hC8;
			14'd4356: ff_rdata <= 8'hCD;
			14'd4357: ff_rdata <= 8'h0F;
			14'd4358: ff_rdata <= 8'h51;
			14'd4359: ff_rdata <= 8'hCD;
			14'd4360: ff_rdata <= 8'h0D;
			14'd4361: ff_rdata <= 8'h51;
			14'd4362: ff_rdata <= 8'hFB;
			14'd4363: ff_rdata <= 8'hB7;
			14'd4364: ff_rdata <= 8'hC9;
			14'd4365: ff_rdata <= 8'hD5;
			14'd4366: ff_rdata <= 8'hC9;
			14'd4367: ff_rdata <= 8'hE5;
			14'd4368: ff_rdata <= 8'hD5;
			14'd4369: ff_rdata <= 8'h21;
			14'd4370: ff_rdata <= 8'h00;
			14'd4371: ff_rdata <= 8'hFD;
			14'd4372: ff_rdata <= 8'h39;
			14'd4373: ff_rdata <= 8'hD2;
			14'd4374: ff_rdata <= 8'h79;
			14'd4375: ff_rdata <= 8'h67;
			14'd4376: ff_rdata <= 8'hED;
			14'd4377: ff_rdata <= 8'h5B;
			14'd4378: ff_rdata <= 8'hC6;
			14'd4379: ff_rdata <= 8'hF6;
			14'd4380: ff_rdata <= 8'hB7;
			14'd4381: ff_rdata <= 8'hED;
			14'd4382: ff_rdata <= 8'h52;
			14'd4383: ff_rdata <= 8'hDA;
			14'd4384: ff_rdata <= 8'h79;
			14'd4385: ff_rdata <= 8'h67;
			14'd4386: ff_rdata <= 8'hD1;
			14'd4387: ff_rdata <= 8'hE1;
			14'd4388: ff_rdata <= 8'hC9;
			14'd4389: ff_rdata <= 8'h00;
			14'd4390: ff_rdata <= 8'h1E;
			14'd4391: ff_rdata <= 8'h23;
			14'd4392: ff_rdata <= 8'h1D;
			14'd4393: ff_rdata <= 8'h1D;
			14'd4394: ff_rdata <= 8'h1D;
			14'd4395: ff_rdata <= 8'h1D;
			14'd4396: ff_rdata <= 8'h1D;
			14'd4397: ff_rdata <= 8'h41;
			14'd4398: ff_rdata <= 8'h1D;
			14'd4399: ff_rdata <= 8'h47;
			14'd4400: ff_rdata <= 8'h57;
			14'd4401: ff_rdata <= 8'h61;
			14'd4402: ff_rdata <= 8'h1D;
			14'd4403: ff_rdata <= 8'h1D;
			14'd4404: ff_rdata <= 8'hF1;
			14'd4405: ff_rdata <= 8'h1D;
			14'd4406: ff_rdata <= 8'h97;
			14'd4407: ff_rdata <= 8'hAE;
			14'd4408: ff_rdata <= 8'hCD;
			14'd4409: ff_rdata <= 8'h1D;
			14'd4410: ff_rdata <= 8'hDF;
			14'd4411: ff_rdata <= 8'h55;
			14'd4412: ff_rdata <= 8'h44;
			14'd4413: ff_rdata <= 8'h52;
			14'd4414: ff_rdata <= 8'h45;
			14'd4415: ff_rdata <= 8'hC7;
			14'd4416: ff_rdata <= 8'h98;
			14'd4417: ff_rdata <= 8'h54;
			14'd4418: ff_rdata <= 8'h50;
			14'd4419: ff_rdata <= 8'h50;
			14'd4420: ff_rdata <= 8'h45;
			14'd4421: ff_rdata <= 8'h4E;
			14'd4422: ff_rdata <= 8'h44;
			14'd4423: ff_rdata <= 8'hFF;
			14'd4424: ff_rdata <= 8'h4D;
			14'd4425: ff_rdata <= 8'hCB;
			14'd4426: ff_rdata <= 8'hB1;
			14'd4427: ff_rdata <= 8'h52;
			14'd4428: ff_rdata <= 8'h50;
			14'd4429: ff_rdata <= 8'h45;
			14'd4430: ff_rdata <= 8'h45;
			14'd4431: ff_rdata <= 8'hCB;
			14'd4432: ff_rdata <= 8'hB1;
			14'd4433: ff_rdata <= 8'h52;
			14'd4434: ff_rdata <= 8'h50;
			14'd4435: ff_rdata <= 8'h4F;
			14'd4436: ff_rdata <= 8'h4B;
			14'd4437: ff_rdata <= 8'hC5;
			14'd4438: ff_rdata <= 8'hB1;
			14'd4439: ff_rdata <= 8'h52;
			14'd4440: ff_rdata <= 8'hFF;
			14'd4441: ff_rdata <= 8'h47;
			14'd4442: ff_rdata <= 8'hCD;
			14'd4443: ff_rdata <= 8'h58;
			14'd4444: ff_rdata <= 8'h54;
			14'd4445: ff_rdata <= 8'hFF;
			14'd4446: ff_rdata <= 8'h4F;
			14'd4447: ff_rdata <= 8'h4E;
			14'd4448: ff_rdata <= 8'h54;
			14'd4449: ff_rdata <= 8'hFF;
			14'd4450: ff_rdata <= 8'h4D;
			14'd4451: ff_rdata <= 8'hCB;
			14'd4452: ff_rdata <= 8'hB1;
			14'd4453: ff_rdata <= 8'h52;
			14'd4454: ff_rdata <= 8'h4F;
			14'd4455: ff_rdata <= 8'h50;
			14'd4456: ff_rdata <= 8'h59;
			14'd4457: ff_rdata <= 8'hFF;
			14'd4458: ff_rdata <= 8'h50;
			14'd4459: ff_rdata <= 8'h43;
			14'd4460: ff_rdata <= 8'hCD;
			14'd4461: ff_rdata <= 8'hB1;
			14'd4462: ff_rdata <= 8'h52;
			14'd4463: ff_rdata <= 8'h4F;
			14'd4464: ff_rdata <= 8'h4E;
			14'd4465: ff_rdata <= 8'h56;
			14'd4466: ff_rdata <= 8'hD0;
			14'd4467: ff_rdata <= 8'hB1;
			14'd4468: ff_rdata <= 8'h52;
			14'd4469: ff_rdata <= 8'h4F;
			14'd4470: ff_rdata <= 8'h4E;
			14'd4471: ff_rdata <= 8'h56;
			14'd4472: ff_rdata <= 8'hC1;
			14'd4473: ff_rdata <= 8'hB1;
			14'd4474: ff_rdata <= 8'h52;
			14'd4475: ff_rdata <= 8'hFF;
			14'd4476: ff_rdata <= 8'h4E;
			14'd4477: ff_rdata <= 8'h4D;
			14'd4478: ff_rdata <= 8'hCB;
			14'd4479: ff_rdata <= 8'hB1;
			14'd4480: ff_rdata <= 8'h52;
			14'd4481: ff_rdata <= 8'hFF;
			14'd4482: ff_rdata <= 8'h45;
			14'd4483: ff_rdata <= 8'h59;
			14'd4484: ff_rdata <= 8'hFF;
			14'd4485: ff_rdata <= 8'h4F;
			14'd4486: ff_rdata <= 8'hCE;
			14'd4487: ff_rdata <= 8'hB1;
			14'd4488: ff_rdata <= 8'h52;
			14'd4489: ff_rdata <= 8'h45;
			14'd4490: ff_rdata <= 8'h59;
			14'd4491: ff_rdata <= 8'hFF;
			14'd4492: ff_rdata <= 8'h4F;
			14'd4493: ff_rdata <= 8'h46;
			14'd4494: ff_rdata <= 8'hC6;
			14'd4495: ff_rdata <= 8'hB1;
			14'd4496: ff_rdata <= 8'h52;
			14'd4497: ff_rdata <= 8'hFF;
			14'd4498: ff_rdata <= 8'h4F;
			14'd4499: ff_rdata <= 8'h41;
			14'd4500: ff_rdata <= 8'h44;
			14'd4501: ff_rdata <= 8'hFF;
			14'd4502: ff_rdata <= 8'h50;
			14'd4503: ff_rdata <= 8'h43;
			14'd4504: ff_rdata <= 8'hCD;
			14'd4505: ff_rdata <= 8'hB1;
			14'd4506: ff_rdata <= 8'h52;
			14'd4507: ff_rdata <= 8'hFF;
			14'd4508: ff_rdata <= 8'h4B;
			14'd4509: ff_rdata <= 8'hFF;
			14'd4510: ff_rdata <= 8'h56;
			14'd4511: ff_rdata <= 8'h4F;
			14'd4512: ff_rdata <= 8'h49;
			14'd4513: ff_rdata <= 8'h43;
			14'd4514: ff_rdata <= 8'hC5;
			14'd4515: ff_rdata <= 8'hB1;
			14'd4516: ff_rdata <= 8'h52;
			14'd4517: ff_rdata <= 8'h4B;
			14'd4518: ff_rdata <= 8'hFF;
			14'd4519: ff_rdata <= 8'h56;
			14'd4520: ff_rdata <= 8'h45;
			14'd4521: ff_rdata <= 8'hCC;
			14'd4522: ff_rdata <= 8'hB1;
			14'd4523: ff_rdata <= 8'h52;
			14'd4524: ff_rdata <= 8'h4B;
			14'd4525: ff_rdata <= 8'hFF;
			14'd4526: ff_rdata <= 8'h56;
			14'd4527: ff_rdata <= 8'h4F;
			14'd4528: ff_rdata <= 8'hCC;
			14'd4529: ff_rdata <= 8'hB1;
			14'd4530: ff_rdata <= 8'h52;
			14'd4531: ff_rdata <= 8'h4B;
			14'd4532: ff_rdata <= 8'hFF;
			14'd4533: ff_rdata <= 8'h54;
			14'd4534: ff_rdata <= 8'h45;
			14'd4535: ff_rdata <= 8'h4D;
			14'd4536: ff_rdata <= 8'h50;
			14'd4537: ff_rdata <= 8'hCF;
			14'd4538: ff_rdata <= 8'hB1;
			14'd4539: ff_rdata <= 8'h52;
			14'd4540: ff_rdata <= 8'h4B;
			14'd4541: ff_rdata <= 8'hFF;
			14'd4542: ff_rdata <= 8'h53;
			14'd4543: ff_rdata <= 8'h54;
			14'd4544: ff_rdata <= 8'h41;
			14'd4545: ff_rdata <= 8'hD4;
			14'd4546: ff_rdata <= 8'hB1;
			14'd4547: ff_rdata <= 8'h52;
			14'd4548: ff_rdata <= 8'h4B;
			14'd4549: ff_rdata <= 8'hFF;
			14'd4550: ff_rdata <= 8'h50;
			14'd4551: ff_rdata <= 8'h43;
			14'd4552: ff_rdata <= 8'hCD;
			14'd4553: ff_rdata <= 8'hB1;
			14'd4554: ff_rdata <= 8'h52;
			14'd4555: ff_rdata <= 8'h55;
			14'd4556: ff_rdata <= 8'h53;
			14'd4557: ff_rdata <= 8'h49;
			14'd4558: ff_rdata <= 8'hC3;
			14'd4559: ff_rdata <= 8'hEC;
			14'd4560: ff_rdata <= 8'h52;
			14'd4561: ff_rdata <= 8'hFF;
			14'd4562: ff_rdata <= 8'h45;
			14'd4563: ff_rdata <= 8'h43;
			14'd4564: ff_rdata <= 8'hFF;
			14'd4565: ff_rdata <= 8'h4D;
			14'd4566: ff_rdata <= 8'hCB;
			14'd4567: ff_rdata <= 8'hB1;
			14'd4568: ff_rdata <= 8'h52;
			14'd4569: ff_rdata <= 8'h45;
			14'd4570: ff_rdata <= 8'h43;
			14'd4571: ff_rdata <= 8'h4D;
			14'd4572: ff_rdata <= 8'h4F;
			14'd4573: ff_rdata <= 8'hC4;
			14'd4574: ff_rdata <= 8'hB1;
			14'd4575: ff_rdata <= 8'h52;
			14'd4576: ff_rdata <= 8'h45;
			14'd4577: ff_rdata <= 8'h43;
			14'd4578: ff_rdata <= 8'hFF;
			14'd4579: ff_rdata <= 8'h50;
			14'd4580: ff_rdata <= 8'h43;
			14'd4581: ff_rdata <= 8'hCD;
			14'd4582: ff_rdata <= 8'hB1;
			14'd4583: ff_rdata <= 8'h52;
			14'd4584: ff_rdata <= 8'hFF;
			14'd4585: ff_rdata <= 8'h54;
			14'd4586: ff_rdata <= 8'h4F;
			14'd4587: ff_rdata <= 8'h50;
			14'd4588: ff_rdata <= 8'hCD;
			14'd4589: ff_rdata <= 8'h8B;
			14'd4590: ff_rdata <= 8'h54;
			14'd4591: ff_rdata <= 8'h45;
			14'd4592: ff_rdata <= 8'h54;
			14'd4593: ff_rdata <= 8'hFF;
			14'd4594: ff_rdata <= 8'h50;
			14'd4595: ff_rdata <= 8'h43;
			14'd4596: ff_rdata <= 8'hCD;
			14'd4597: ff_rdata <= 8'hB1;
			14'd4598: ff_rdata <= 8'h52;
			14'd4599: ff_rdata <= 8'h41;
			14'd4600: ff_rdata <= 8'h56;
			14'd4601: ff_rdata <= 8'h45;
			14'd4602: ff_rdata <= 8'hFF;
			14'd4603: ff_rdata <= 8'h50;
			14'd4604: ff_rdata <= 8'h43;
			14'd4605: ff_rdata <= 8'hCD;
			14'd4606: ff_rdata <= 8'hB1;
			14'd4607: ff_rdata <= 8'h52;
			14'd4608: ff_rdata <= 8'h59;
			14'd4609: ff_rdata <= 8'h4E;
			14'd4610: ff_rdata <= 8'h54;
			14'd4611: ff_rdata <= 8'h48;
			14'd4612: ff_rdata <= 8'hC5;
			14'd4613: ff_rdata <= 8'hB1;
			14'd4614: ff_rdata <= 8'h52;
			14'd4615: ff_rdata <= 8'hFF;
			14'd4616: ff_rdata <= 8'h52;
			14'd4617: ff_rdata <= 8'h41;
			14'd4618: ff_rdata <= 8'h4E;
			14'd4619: ff_rdata <= 8'h53;
			14'd4620: ff_rdata <= 8'h50;
			14'd4621: ff_rdata <= 8'h4F;
			14'd4622: ff_rdata <= 8'h53;
			14'd4623: ff_rdata <= 8'hC5;
			14'd4624: ff_rdata <= 8'h35;
			14'd4625: ff_rdata <= 8'h55;
			14'd4626: ff_rdata <= 8'h45;
			14'd4627: ff_rdata <= 8'h4D;
			14'd4628: ff_rdata <= 8'h50;
			14'd4629: ff_rdata <= 8'h45;
			14'd4630: ff_rdata <= 8'hD2;
			14'd4631: ff_rdata <= 8'h41;
			14'd4632: ff_rdata <= 8'h55;
			14'd4633: ff_rdata <= 8'hFF;
			14'd4634: ff_rdata <= 8'h4F;
			14'd4635: ff_rdata <= 8'h49;
			14'd4636: ff_rdata <= 8'h43;
			14'd4637: ff_rdata <= 8'hC5;
			14'd4638: ff_rdata <= 8'hEE;
			14'd4639: ff_rdata <= 8'h55;
			14'd4640: ff_rdata <= 8'h4F;
			14'd4641: ff_rdata <= 8'h49;
			14'd4642: ff_rdata <= 8'h43;
			14'd4643: ff_rdata <= 8'h45;
			14'd4644: ff_rdata <= 8'hFF;
			14'd4645: ff_rdata <= 8'h43;
			14'd4646: ff_rdata <= 8'h4F;
			14'd4647: ff_rdata <= 8'h50;
			14'd4648: ff_rdata <= 8'hD9;
			14'd4649: ff_rdata <= 8'h7E;
			14'd4650: ff_rdata <= 8'h56;
			14'd4651: ff_rdata <= 8'hFF;
			14'd4652: ff_rdata <= 8'h4C;
			14'd4653: ff_rdata <= 8'h41;
			14'd4654: ff_rdata <= 8'hD9;
			14'd4655: ff_rdata <= 8'h46;
			14'd4656: ff_rdata <= 8'h57;
			14'd4657: ff_rdata <= 8'h4C;
			14'd4658: ff_rdata <= 8'h41;
			14'd4659: ff_rdata <= 8'h59;
			14'd4660: ff_rdata <= 8'hFF;
			14'd4661: ff_rdata <= 8'h50;
			14'd4662: ff_rdata <= 8'h43;
			14'd4663: ff_rdata <= 8'hCD;
			14'd4664: ff_rdata <= 8'hB1;
			14'd4665: ff_rdata <= 8'h52;
			14'd4666: ff_rdata <= 8'h43;
			14'd4667: ff_rdata <= 8'h4D;
			14'd4668: ff_rdata <= 8'hFF;
			14'd4669: ff_rdata <= 8'h46;
			14'd4670: ff_rdata <= 8'h52;
			14'd4671: ff_rdata <= 8'h45;
			14'd4672: ff_rdata <= 8'hD1;
			14'd4673: ff_rdata <= 8'hB1;
			14'd4674: ff_rdata <= 8'h52;
			14'd4675: ff_rdata <= 8'h43;
			14'd4676: ff_rdata <= 8'h4D;
			14'd4677: ff_rdata <= 8'hFF;
			14'd4678: ff_rdata <= 8'h56;
			14'd4679: ff_rdata <= 8'h4F;
			14'd4680: ff_rdata <= 8'hCC;
			14'd4681: ff_rdata <= 8'hB1;
			14'd4682: ff_rdata <= 8'h52;
			14'd4683: ff_rdata <= 8'h4C;
			14'd4684: ff_rdata <= 8'h41;
			14'd4685: ff_rdata <= 8'h59;
			14'd4686: ff_rdata <= 8'hFF;
			14'd4687: ff_rdata <= 8'h4D;
			14'd4688: ff_rdata <= 8'hCB;
			14'd4689: ff_rdata <= 8'hB1;
			14'd4690: ff_rdata <= 8'h52;
			14'd4691: ff_rdata <= 8'h49;
			14'd4692: ff_rdata <= 8'h54;
			14'd4693: ff_rdata <= 8'h43;
			14'd4694: ff_rdata <= 8'hC8;
			14'd4695: ff_rdata <= 8'h29;
			14'd4696: ff_rdata <= 8'h55;
			14'd4697: ff_rdata <= 8'hFF;
			14'd4698: ff_rdata <= 8'h7E;
			14'd4699: ff_rdata <= 8'hD6;
			14'd4700: ff_rdata <= 8'h41;
			14'd4701: ff_rdata <= 8'hD8;
			14'd4702: ff_rdata <= 8'hFE;
			14'd4703: ff_rdata <= 8'h16;
			14'd4704: ff_rdata <= 8'h3F;
			14'd4705: ff_rdata <= 8'hD8;
			14'd4706: ff_rdata <= 8'h23;
			14'd4707: ff_rdata <= 8'hE5;
			14'd4708: ff_rdata <= 8'h21;
			14'd4709: ff_rdata <= 8'h25;
			14'd4710: ff_rdata <= 8'h51;
			14'd4711: ff_rdata <= 8'hCD;
			14'd4712: ff_rdata <= 8'h86;
			14'd4713: ff_rdata <= 8'h54;
			14'd4714: ff_rdata <= 8'h7E;
			14'd4715: ff_rdata <= 8'h21;
			14'd4716: ff_rdata <= 8'h3B;
			14'd4717: ff_rdata <= 8'h51;
			14'd4718: ff_rdata <= 8'hCD;
			14'd4719: ff_rdata <= 8'h86;
			14'd4720: ff_rdata <= 8'h54;
			14'd4721: ff_rdata <= 8'hEB;
			14'd4722: ff_rdata <= 8'hE1;
			14'd4723: ff_rdata <= 8'hE5;
			14'd4724: ff_rdata <= 8'h1A;
			14'd4725: ff_rdata <= 8'h3C;
			14'd4726: ff_rdata <= 8'h28;
			14'd4727: ff_rdata <= 8'h0B;
			14'd4728: ff_rdata <= 8'hCD;
			14'd4729: ff_rdata <= 8'h86;
			14'd4730: ff_rdata <= 8'h52;
			14'd4731: ff_rdata <= 8'hE1;
			14'd4732: ff_rdata <= 8'h20;
			14'd4733: ff_rdata <= 8'hF5;
			14'd4734: ff_rdata <= 8'hEB;
			14'd4735: ff_rdata <= 8'h5E;
			14'd4736: ff_rdata <= 8'h23;
			14'd4737: ff_rdata <= 8'h56;
			14'd4738: ff_rdata <= 8'hC9;
			14'd4739: ff_rdata <= 8'h37;
			14'd4740: ff_rdata <= 8'hE1;
			14'd4741: ff_rdata <= 8'hC9;
			14'd4742: ff_rdata <= 8'h1A;
			14'd4743: ff_rdata <= 8'h47;
			14'd4744: ff_rdata <= 8'hE6;
			14'd4745: ff_rdata <= 8'h7F;
			14'd4746: ff_rdata <= 8'hBE;
			14'd4747: ff_rdata <= 8'h13;
			14'd4748: ff_rdata <= 8'h23;
			14'd4749: ff_rdata <= 8'h20;
			14'd4750: ff_rdata <= 8'h08;
			14'd4751: ff_rdata <= 8'h78;
			14'd4752: ff_rdata <= 8'hB7;
			14'd4753: ff_rdata <= 8'hF2;
			14'd4754: ff_rdata <= 8'h86;
			14'd4755: ff_rdata <= 8'h52;
			14'd4756: ff_rdata <= 8'h7E;
			14'd4757: ff_rdata <= 8'hB7;
			14'd4758: ff_rdata <= 8'hC8;
			14'd4759: ff_rdata <= 8'h04;
			14'd4760: ff_rdata <= 8'h20;
			14'd4761: ff_rdata <= 8'h0A;
			14'd4762: ff_rdata <= 8'h2B;
			14'd4763: ff_rdata <= 8'h7E;
			14'd4764: ff_rdata <= 8'hFE;
			14'd4765: ff_rdata <= 8'h20;
			14'd4766: ff_rdata <= 8'h23;
			14'd4767: ff_rdata <= 8'h28;
			14'd4768: ff_rdata <= 8'hFA;
			14'd4769: ff_rdata <= 8'h2B;
			14'd4770: ff_rdata <= 8'h18;
			14'd4771: ff_rdata <= 8'hE2;
			14'd4772: ff_rdata <= 8'h1B;
			14'd4773: ff_rdata <= 8'h1A;
			14'd4774: ff_rdata <= 8'h13;
			14'd4775: ff_rdata <= 8'h3C;
			14'd4776: ff_rdata <= 8'h28;
			14'd4777: ff_rdata <= 8'hFB;
			14'd4778: ff_rdata <= 8'h3D;
			14'd4779: ff_rdata <= 8'hF2;
			14'd4780: ff_rdata <= 8'hA5;
			14'd4781: ff_rdata <= 8'h52;
			14'd4782: ff_rdata <= 8'h13;
			14'd4783: ff_rdata <= 8'h13;
			14'd4784: ff_rdata <= 8'hC9;
			14'd4785: ff_rdata <= 8'hC3;
			14'd4786: ff_rdata <= 8'h70;
			14'd4787: ff_rdata <= 8'h67;
			14'd4788: ff_rdata <= 8'hCD;
			14'd4789: ff_rdata <= 8'hE4;
			14'd4790: ff_rdata <= 8'h55;
			14'd4791: ff_rdata <= 8'hC3;
			14'd4792: ff_rdata <= 8'hC1;
			14'd4793: ff_rdata <= 8'h67;
			14'd4794: ff_rdata <= 8'hCD;
			14'd4795: ff_rdata <= 8'hE7;
			14'd4796: ff_rdata <= 8'h54;
			14'd4797: ff_rdata <= 8'hC2;
			14'd4798: ff_rdata <= 8'h6D;
			14'd4799: ff_rdata <= 8'h67;
			14'd4800: ff_rdata <= 8'hC9;
			14'd4801: ff_rdata <= 8'hC5;
			14'd4802: ff_rdata <= 8'hCD;
			14'd4803: ff_rdata <= 8'hB4;
			14'd4804: ff_rdata <= 8'h52;
			14'd4805: ff_rdata <= 8'h18;
			14'd4806: ff_rdata <= 8'h13;
			14'd4807: ff_rdata <= 8'hC5;
			14'd4808: ff_rdata <= 8'hCD;
			14'd4809: ff_rdata <= 8'hE4;
			14'd4810: ff_rdata <= 8'h55;
			14'd4811: ff_rdata <= 8'h18;
			14'd4812: ff_rdata <= 8'h0A;
			14'd4813: ff_rdata <= 8'hCD;
			14'd4814: ff_rdata <= 8'hE4;
			14'd4815: ff_rdata <= 8'h55;
			14'd4816: ff_rdata <= 8'hCD;
			14'd4817: ff_rdata <= 8'hBB;
			14'd4818: ff_rdata <= 8'h67;
			14'd4819: ff_rdata <= 8'hD5;
			14'd4820: ff_rdata <= 8'hCD;
			14'd4821: ff_rdata <= 8'hDF;
			14'd4822: ff_rdata <= 8'h55;
			14'd4823: ff_rdata <= 8'hCD;
			14'd4824: ff_rdata <= 8'hBB;
			14'd4825: ff_rdata <= 8'h67;
			14'd4826: ff_rdata <= 8'hCD;
			14'd4827: ff_rdata <= 8'hE9;
			14'd4828: ff_rdata <= 8'h55;
			14'd4829: ff_rdata <= 8'hC1;
			14'd4830: ff_rdata <= 8'h7B;
			14'd4831: ff_rdata <= 8'hC9;
			14'd4832: ff_rdata <= 8'h03;
			14'd4833: ff_rdata <= 8'h01;
			14'd4834: ff_rdata <= 8'h00;
			14'd4835: ff_rdata <= 8'h01;
			14'd4836: ff_rdata <= 8'h01;
			14'd4837: ff_rdata <= 8'h01;
			14'd4838: ff_rdata <= 8'h00;
			14'd4839: ff_rdata <= 8'h00;
			14'd4840: ff_rdata <= 8'h00;
			14'd4841: ff_rdata <= 8'h00;
			14'd4842: ff_rdata <= 8'h00;
			14'd4843: ff_rdata <= 8'h00;
			14'd4844: ff_rdata <= 8'hE5;
			14'd4845: ff_rdata <= 8'hCD;
			14'd4846: ff_rdata <= 8'hC6;
			14'd4847: ff_rdata <= 8'h50;
			14'd4848: ff_rdata <= 8'hCC;
			14'd4849: ff_rdata <= 8'h09;
			14'd4850: ff_rdata <= 8'h50;
			14'd4851: ff_rdata <= 8'h21;
			14'd4852: ff_rdata <= 8'hE0;
			14'd4853: ff_rdata <= 8'h52;
			14'd4854: ff_rdata <= 8'h11;
			14'd4855: ff_rdata <= 8'h5E;
			14'd4856: ff_rdata <= 8'hF5;
			14'd4857: ff_rdata <= 8'h01;
			14'd4858: ff_rdata <= 8'h0C;
			14'd4859: ff_rdata <= 8'h00;
			14'd4860: ff_rdata <= 8'hED;
			14'd4861: ff_rdata <= 8'hB0;
			14'd4862: ff_rdata <= 8'hE1;
			14'd4863: ff_rdata <= 8'hCD;
			14'd4864: ff_rdata <= 8'hE7;
			14'd4865: ff_rdata <= 8'h54;
			14'd4866: ff_rdata <= 8'h28;
			14'd4867: ff_rdata <= 8'h6B;
			14'd4868: ff_rdata <= 8'hE5;
			14'd4869: ff_rdata <= 8'h21;
			14'd4870: ff_rdata <= 8'h5E;
			14'd4871: ff_rdata <= 8'hF5;
			14'd4872: ff_rdata <= 8'h11;
			14'd4873: ff_rdata <= 8'h5F;
			14'd4874: ff_rdata <= 8'hF5;
			14'd4875: ff_rdata <= 8'h01;
			14'd4876: ff_rdata <= 8'h0B;
			14'd4877: ff_rdata <= 8'h00;
			14'd4878: ff_rdata <= 8'h36;
			14'd4879: ff_rdata <= 8'h00;
			14'd4880: ff_rdata <= 8'hED;
			14'd4881: ff_rdata <= 8'hB0;
			14'd4882: ff_rdata <= 8'hE1;
			14'd4883: ff_rdata <= 8'hCD;
			14'd4884: ff_rdata <= 8'hE4;
			14'd4885: ff_rdata <= 8'h55;
			14'd4886: ff_rdata <= 8'hFE;
			14'd4887: ff_rdata <= 8'h2C;
			14'd4888: ff_rdata <= 8'h28;
			14'd4889: ff_rdata <= 8'h10;
			14'd4890: ff_rdata <= 8'hCD;
			14'd4891: ff_rdata <= 8'hC1;
			14'd4892: ff_rdata <= 8'h67;
			14'd4893: ff_rdata <= 8'hFE;
			14'd4894: ff_rdata <= 8'h02;
			14'd4895: ff_rdata <= 8'hD2;
			14'd4896: ff_rdata <= 8'h70;
			14'd4897: ff_rdata <= 8'h67;
			14'd4898: ff_rdata <= 8'h32;
			14'd4899: ff_rdata <= 8'h5F;
			14'd4900: ff_rdata <= 8'hF5;
			14'd4901: ff_rdata <= 8'h7E;
			14'd4902: ff_rdata <= 8'hFE;
			14'd4903: ff_rdata <= 8'h29;
			14'd4904: ff_rdata <= 8'h28;
			14'd4905: ff_rdata <= 8'h3F;
			14'd4906: ff_rdata <= 8'hCD;
			14'd4907: ff_rdata <= 8'hDF;
			14'd4908: ff_rdata <= 8'h55;
			14'd4909: ff_rdata <= 8'hFE;
			14'd4910: ff_rdata <= 8'h2C;
			14'd4911: ff_rdata <= 8'h28;
			14'd4912: ff_rdata <= 8'h0E;
			14'd4913: ff_rdata <= 8'hCD;
			14'd4914: ff_rdata <= 8'hC1;
			14'd4915: ff_rdata <= 8'h67;
			14'd4916: ff_rdata <= 8'hB7;
			14'd4917: ff_rdata <= 8'h20;
			14'd4918: ff_rdata <= 8'h1E;
			14'd4919: ff_rdata <= 8'h32;
			14'd4920: ff_rdata <= 8'h60;
			14'd4921: ff_rdata <= 8'hF5;
			14'd4922: ff_rdata <= 8'h7E;
			14'd4923: ff_rdata <= 8'hFE;
			14'd4924: ff_rdata <= 8'h29;
			14'd4925: ff_rdata <= 8'h28;
			14'd4926: ff_rdata <= 8'h2A;
			14'd4927: ff_rdata <= 8'h06;
			14'd4928: ff_rdata <= 8'h09;
			14'd4929: ff_rdata <= 8'hE5;
			14'd4930: ff_rdata <= 8'h21;
			14'd4931: ff_rdata <= 8'h61;
			14'd4932: ff_rdata <= 8'hF5;
			14'd4933: ff_rdata <= 8'hE3;
			14'd4934: ff_rdata <= 8'h0E;
			14'd4935: ff_rdata <= 8'h00;
			14'd4936: ff_rdata <= 8'hCD;
			14'd4937: ff_rdata <= 8'hDF;
			14'd4938: ff_rdata <= 8'h55;
			14'd4939: ff_rdata <= 8'hC5;
			14'd4940: ff_rdata <= 8'hCD;
			14'd4941: ff_rdata <= 8'hC1;
			14'd4942: ff_rdata <= 8'h67;
			14'd4943: ff_rdata <= 8'hC1;
			14'd4944: ff_rdata <= 8'hB7;
			14'd4945: ff_rdata <= 8'h28;
			14'd4946: ff_rdata <= 8'h02;
			14'd4947: ff_rdata <= 8'hFE;
			14'd4948: ff_rdata <= 8'h0A;
			14'd4949: ff_rdata <= 8'hD2;
			14'd4950: ff_rdata <= 8'h70;
			14'd4951: ff_rdata <= 8'h67;
			14'd4952: ff_rdata <= 8'hE3;
			14'd4953: ff_rdata <= 8'h77;
			14'd4954: ff_rdata <= 8'h23;
			14'd4955: ff_rdata <= 8'h0C;
			14'd4956: ff_rdata <= 8'hE3;
			14'd4957: ff_rdata <= 8'h7E;
			14'd4958: ff_rdata <= 8'hFE;
			14'd4959: ff_rdata <= 8'h29;
			14'd4960: ff_rdata <= 8'h28;
			14'd4961: ff_rdata <= 8'h02;
			14'd4962: ff_rdata <= 8'h10;
			14'd4963: ff_rdata <= 8'hE4;
			14'd4964: ff_rdata <= 8'h79;
			14'd4965: ff_rdata <= 8'h32;
			14'd4966: ff_rdata <= 8'h5E;
			14'd4967: ff_rdata <= 8'hF5;
			14'd4968: ff_rdata <= 8'hC1;
			14'd4969: ff_rdata <= 8'hCD;
			14'd4970: ff_rdata <= 8'hE9;
			14'd4971: ff_rdata <= 8'h55;
			14'd4972: ff_rdata <= 8'hC2;
			14'd4973: ff_rdata <= 8'h6D;
			14'd4974: ff_rdata <= 8'h67;
			14'd4975: ff_rdata <= 8'hE5;
			14'd4976: ff_rdata <= 8'h21;
			14'd4977: ff_rdata <= 8'h5F;
			14'd4978: ff_rdata <= 8'hF5;
			14'd4979: ff_rdata <= 8'h7E;
			14'd4980: ff_rdata <= 8'hE6;
			14'd4981: ff_rdata <= 8'h01;
			14'd4982: ff_rdata <= 8'h57;
			14'd4983: ff_rdata <= 8'h87;
			14'd4984: ff_rdata <= 8'h82;
			14'd4985: ff_rdata <= 8'h23;
			14'd4986: ff_rdata <= 8'h86;
			14'd4987: ff_rdata <= 8'h23;
			14'd4988: ff_rdata <= 8'h57;
			14'd4989: ff_rdata <= 8'h3A;
			14'd4990: ff_rdata <= 8'h5E;
			14'd4991: ff_rdata <= 8'hF5;
			14'd4992: ff_rdata <= 8'h47;
			14'd4993: ff_rdata <= 8'hB7;
			14'd4994: ff_rdata <= 8'h28;
			14'd4995: ff_rdata <= 8'h05;
			14'd4996: ff_rdata <= 8'hAF;
			14'd4997: ff_rdata <= 8'h86;
			14'd4998: ff_rdata <= 8'h23;
			14'd4999: ff_rdata <= 8'h10;
			14'd5000: ff_rdata <= 8'hFC;
			14'd5001: ff_rdata <= 8'h82;
			14'd5002: ff_rdata <= 8'hFE;
			14'd5003: ff_rdata <= 8'h0A;
			14'd5004: ff_rdata <= 8'h30;
			14'd5005: ff_rdata <= 8'hC7;
			14'd5006: ff_rdata <= 8'hCD;
			14'd5007: ff_rdata <= 8'hCD;
			14'd5008: ff_rdata <= 8'h67;
			14'd5009: ff_rdata <= 8'h2A;
			14'd5010: ff_rdata <= 8'h4A;
			14'd5011: ff_rdata <= 8'hFC;
			14'd5012: ff_rdata <= 8'hCD;
			14'd5013: ff_rdata <= 8'hC6;
			14'd5014: ff_rdata <= 8'h50;
			14'd5015: ff_rdata <= 8'h20;
			14'd5016: ff_rdata <= 8'h16;
			14'd5017: ff_rdata <= 8'h11;
			14'd5018: ff_rdata <= 8'h27;
			14'd5019: ff_rdata <= 8'h03;
			14'd5020: ff_rdata <= 8'hA7;
			14'd5021: ff_rdata <= 8'hED;
			14'd5022: ff_rdata <= 8'h52;
			14'd5023: ff_rdata <= 8'h22;
			14'd5024: ff_rdata <= 8'h4A;
			14'd5025: ff_rdata <= 8'hFC;
			14'd5026: ff_rdata <= 8'h22;
			14'd5027: ff_rdata <= 8'h7D;
			14'd5028: ff_rdata <= 8'hF9;
			14'd5029: ff_rdata <= 8'h3A;
			14'd5030: ff_rdata <= 8'hA7;
			14'd5031: ff_rdata <= 8'hFF;
			14'd5032: ff_rdata <= 8'hFE;
			14'd5033: ff_rdata <= 8'hC9;
			14'd5034: ff_rdata <= 8'h28;
			14'd5035: ff_rdata <= 8'h03;
			14'd5036: ff_rdata <= 8'h22;
			14'd5037: ff_rdata <= 8'h49;
			14'd5038: ff_rdata <= 8'hF3;
			14'd5039: ff_rdata <= 8'hD1;
			14'd5040: ff_rdata <= 8'hF9;
			14'd5041: ff_rdata <= 8'hD5;
			14'd5042: ff_rdata <= 8'hCD;
			14'd5043: ff_rdata <= 8'h07;
			14'd5044: ff_rdata <= 8'h54;
			14'd5045: ff_rdata <= 8'h2A;
			14'd5046: ff_rdata <= 8'h1C;
			14'd5047: ff_rdata <= 8'hF4;
			14'd5048: ff_rdata <= 8'h22;
			14'd5049: ff_rdata <= 8'hBE;
			14'd5050: ff_rdata <= 8'hF6;
			14'd5051: ff_rdata <= 8'h21;
			14'd5052: ff_rdata <= 8'hEC;
			14'd5053: ff_rdata <= 8'h53;
			14'd5054: ff_rdata <= 8'h11;
			14'd5055: ff_rdata <= 8'h06;
			14'd5056: ff_rdata <= 8'hF8;
			14'd5057: ff_rdata <= 8'h01;
			14'd5058: ff_rdata <= 8'h1B;
			14'd5059: ff_rdata <= 8'h00;
			14'd5060: ff_rdata <= 8'hED;
			14'd5061: ff_rdata <= 8'hB0;
			14'd5062: ff_rdata <= 8'h3A;
			14'd5063: ff_rdata <= 8'h5F;
			14'd5064: ff_rdata <= 8'hF8;
			14'd5065: ff_rdata <= 8'h32;
			14'd5066: ff_rdata <= 8'h0B;
			14'd5067: ff_rdata <= 8'hF8;
			14'd5068: ff_rdata <= 8'hE1;
			14'd5069: ff_rdata <= 8'h7D;
			14'd5070: ff_rdata <= 8'h32;
			14'd5071: ff_rdata <= 8'h13;
			14'd5072: ff_rdata <= 8'hF8;
			14'd5073: ff_rdata <= 8'h7C;
			14'd5074: ff_rdata <= 8'h32;
			14'd5075: ff_rdata <= 8'h1B;
			14'd5076: ff_rdata <= 8'hF8;
			14'd5077: ff_rdata <= 8'hAF;
			14'd5078: ff_rdata <= 8'h32;
			14'd5079: ff_rdata <= 8'h5F;
			14'd5080: ff_rdata <= 8'hF8;
			14'd5081: ff_rdata <= 8'h21;
			14'd5082: ff_rdata <= 8'h5E;
			14'd5083: ff_rdata <= 8'hF5;
			14'd5084: ff_rdata <= 8'h22;
			14'd5085: ff_rdata <= 8'h60;
			14'd5086: ff_rdata <= 8'hF8;
			14'd5087: ff_rdata <= 8'h21;
			14'd5088: ff_rdata <= 8'h60;
			14'd5089: ff_rdata <= 8'hF5;
			14'd5090: ff_rdata <= 8'h22;
			14'd5091: ff_rdata <= 8'h5E;
			14'd5092: ff_rdata <= 8'hF5;
			14'd5093: ff_rdata <= 8'h77;
			14'd5094: ff_rdata <= 8'h21;
			14'd5095: ff_rdata <= 8'h06;
			14'd5096: ff_rdata <= 8'hF8;
			14'd5097: ff_rdata <= 8'hC3;
			14'd5098: ff_rdata <= 8'hC7;
			14'd5099: ff_rdata <= 8'h67;
			14'd5100: ff_rdata <= 8'h3A;
			14'd5101: ff_rdata <= 8'hCD;
			14'd5102: ff_rdata <= 8'hB7;
			14'd5103: ff_rdata <= 8'hEF;
			14'd5104: ff_rdata <= 8'h0F;
			14'd5105: ff_rdata <= 8'h00;
			14'd5106: ff_rdata <= 8'h3A;
			14'd5107: ff_rdata <= 8'h98;
			14'd5108: ff_rdata <= 8'h0C;
			14'd5109: ff_rdata <= 8'hC0;
			14'd5110: ff_rdata <= 8'hF6;
			14'd5111: ff_rdata <= 8'h2C;
			14'd5112: ff_rdata <= 8'h0F;
			14'd5113: ff_rdata <= 8'h00;
			14'd5114: ff_rdata <= 8'h3A;
			14'd5115: ff_rdata <= 8'h98;
			14'd5116: ff_rdata <= 8'h0C;
			14'd5117: ff_rdata <= 8'hC1;
			14'd5118: ff_rdata <= 8'hF6;
			14'd5119: ff_rdata <= 8'h2C;
			14'd5120: ff_rdata <= 8'h0F;
			14'd5121: ff_rdata <= 8'h00;
			14'd5122: ff_rdata <= 8'h3A;
			14'd5123: ff_rdata <= 8'h99;
			14'd5124: ff_rdata <= 8'h00;
			14'd5125: ff_rdata <= 8'h00;
			14'd5126: ff_rdata <= 8'h00;
			14'd5127: ff_rdata <= 8'hF3;
			14'd5128: ff_rdata <= 8'h21;
			14'd5129: ff_rdata <= 8'h5E;
			14'd5130: ff_rdata <= 8'hF5;
			14'd5131: ff_rdata <= 8'h7E;
			14'd5132: ff_rdata <= 8'h32;
			14'd5133: ff_rdata <= 8'h84;
			14'd5134: ff_rdata <= 8'hF9;
			14'd5135: ff_rdata <= 8'h23;
			14'd5136: ff_rdata <= 8'hE5;
			14'd5137: ff_rdata <= 8'h23;
			14'd5138: ff_rdata <= 8'h23;
			14'd5139: ff_rdata <= 8'h11;
			14'd5140: ff_rdata <= 8'h85;
			14'd5141: ff_rdata <= 8'hF9;
			14'd5142: ff_rdata <= 8'h01;
			14'd5143: ff_rdata <= 8'h09;
			14'd5144: ff_rdata <= 8'h00;
			14'd5145: ff_rdata <= 8'hED;
			14'd5146: ff_rdata <= 8'hB0;
			14'd5147: ff_rdata <= 8'hE1;
			14'd5148: ff_rdata <= 8'h46;
			14'd5149: ff_rdata <= 8'h23;
			14'd5150: ff_rdata <= 8'h7E;
			14'd5151: ff_rdata <= 8'h21;
			14'd5152: ff_rdata <= 8'h00;
			14'd5153: ff_rdata <= 8'h00;
			14'd5154: ff_rdata <= 8'hB7;
			14'd5155: ff_rdata <= 8'h28;
			14'd5156: ff_rdata <= 8'h08;
			14'd5157: ff_rdata <= 8'h37;
			14'd5158: ff_rdata <= 8'hCB;
			14'd5159: ff_rdata <= 8'h1C;
			14'd5160: ff_rdata <= 8'hCB;
			14'd5161: ff_rdata <= 8'h1D;
			14'd5162: ff_rdata <= 8'h3D;
			14'd5163: ff_rdata <= 8'h18;
			14'd5164: ff_rdata <= 8'hF6;
			14'd5165: ff_rdata <= 8'h29;
			14'd5166: ff_rdata <= 8'hCB;
			14'd5167: ff_rdata <= 8'h17;
			14'd5168: ff_rdata <= 8'h6C;
			14'd5169: ff_rdata <= 8'h67;
			14'd5170: ff_rdata <= 8'h78;
			14'd5171: ff_rdata <= 8'h32;
			14'd5172: ff_rdata <= 8'h8E;
			14'd5173: ff_rdata <= 8'hF9;
			14'd5174: ff_rdata <= 8'hE6;
			14'd5175: ff_rdata <= 8'h01;
			14'd5176: ff_rdata <= 8'h28;
			14'd5177: ff_rdata <= 8'h0C;
			14'd5178: ff_rdata <= 8'hCB;
			14'd5179: ff_rdata <= 8'h3C;
			14'd5180: ff_rdata <= 8'hCB;
			14'd5181: ff_rdata <= 8'h1D;
			14'd5182: ff_rdata <= 8'hCB;
			14'd5183: ff_rdata <= 8'h3C;
			14'd5184: ff_rdata <= 8'hCB;
			14'd5185: ff_rdata <= 8'h1D;
			14'd5186: ff_rdata <= 8'hCB;
			14'd5187: ff_rdata <= 8'h3C;
			14'd5188: ff_rdata <= 8'hCB;
			14'd5189: ff_rdata <= 8'h1D;
			14'd5190: ff_rdata <= 8'hEB;
			14'd5191: ff_rdata <= 8'hD5;
			14'd5192: ff_rdata <= 8'hCD;
			14'd5193: ff_rdata <= 8'h89;
			14'd5194: ff_rdata <= 8'h64;
			14'd5195: ff_rdata <= 8'hCD;
			14'd5196: ff_rdata <= 8'hEE;
			14'd5197: ff_rdata <= 8'h64;
			14'd5198: ff_rdata <= 8'hCD;
			14'd5199: ff_rdata <= 8'h7F;
			14'd5200: ff_rdata <= 8'h50;
			14'd5201: ff_rdata <= 8'hD1;
			14'd5202: ff_rdata <= 8'hCD;
			14'd5203: ff_rdata <= 8'h84;
			14'd5204: ff_rdata <= 8'h55;
			14'd5205: ff_rdata <= 8'hC3;
			14'd5206: ff_rdata <= 8'h56;
			14'd5207: ff_rdata <= 8'h65;
			14'd5208: ff_rdata <= 8'hCD;
			14'd5209: ff_rdata <= 8'hC1;
			14'd5210: ff_rdata <= 8'h52;
			14'd5211: ff_rdata <= 8'hFE;
			14'd5212: ff_rdata <= 8'h02;
			14'd5213: ff_rdata <= 8'hD2;
			14'd5214: ff_rdata <= 8'h70;
			14'd5215: ff_rdata <= 8'h67;
			14'd5216: ff_rdata <= 8'h3D;
			14'd5217: ff_rdata <= 8'h32;
			14'd5218: ff_rdata <= 8'h98;
			14'd5219: ff_rdata <= 8'hF9;
			14'd5220: ff_rdata <= 8'hC9;
			14'd5221: ff_rdata <= 8'hCD;
			14'd5222: ff_rdata <= 8'hE4;
			14'd5223: ff_rdata <= 8'h55;
			14'd5224: ff_rdata <= 8'hCD;
			14'd5225: ff_rdata <= 8'hBB;
			14'd5226: ff_rdata <= 8'h67;
			14'd5227: ff_rdata <= 8'h7E;
			14'd5228: ff_rdata <= 8'hFE;
			14'd5229: ff_rdata <= 8'h29;
			14'd5230: ff_rdata <= 8'hD5;
			14'd5231: ff_rdata <= 8'h28;
			14'd5232: ff_rdata <= 8'h06;
			14'd5233: ff_rdata <= 8'hCD;
			14'd5234: ff_rdata <= 8'hDF;
			14'd5235: ff_rdata <= 8'h55;
			14'd5236: ff_rdata <= 8'hCD;
			14'd5237: ff_rdata <= 8'hBB;
			14'd5238: ff_rdata <= 8'h67;
			14'd5239: ff_rdata <= 8'hCD;
			14'd5240: ff_rdata <= 8'hE9;
			14'd5241: ff_rdata <= 8'h55;
			14'd5242: ff_rdata <= 8'hC1;
			14'd5243: ff_rdata <= 8'h7B;
			14'd5244: ff_rdata <= 8'hC9;
			14'd5245: ff_rdata <= 8'h7A;
			14'd5246: ff_rdata <= 8'hA7;
			14'd5247: ff_rdata <= 8'h37;
			14'd5248: ff_rdata <= 8'hC0;
			14'd5249: ff_rdata <= 8'h7B;
			14'd5250: ff_rdata <= 8'hFE;
			14'd5251: ff_rdata <= 8'h40;
			14'd5252: ff_rdata <= 8'h3F;
			14'd5253: ff_rdata <= 8'hC9;
			14'd5254: ff_rdata <= 8'h85;
			14'd5255: ff_rdata <= 8'h6F;
			14'd5256: ff_rdata <= 8'hD0;
			14'd5257: ff_rdata <= 8'h24;
			14'd5258: ff_rdata <= 8'hC9;
			14'd5259: ff_rdata <= 8'hCD;
			14'd5260: ff_rdata <= 8'hE7;
			14'd5261: ff_rdata <= 8'h54;
			14'd5262: ff_rdata <= 8'hC2;
			14'd5263: ff_rdata <= 8'h6D;
			14'd5264: ff_rdata <= 8'h67;
			14'd5265: ff_rdata <= 8'hE5;
			14'd5266: ff_rdata <= 8'hCD;
			14'd5267: ff_rdata <= 8'h8D;
			14'd5268: ff_rdata <= 8'h65;
			14'd5269: ff_rdata <= 8'hE1;
			14'd5270: ff_rdata <= 8'hB7;
			14'd5271: ff_rdata <= 8'hC9;
			14'd5272: ff_rdata <= 8'hCD;
			14'd5273: ff_rdata <= 8'hE4;
			14'd5274: ff_rdata <= 8'h55;
			14'd5275: ff_rdata <= 8'hCD;
			14'd5276: ff_rdata <= 8'hC1;
			14'd5277: ff_rdata <= 8'h67;
			14'd5278: ff_rdata <= 8'hD5;
			14'd5279: ff_rdata <= 8'hCD;
			14'd5280: ff_rdata <= 8'hDF;
			14'd5281: ff_rdata <= 8'h55;
			14'd5282: ff_rdata <= 8'hCD;
			14'd5283: ff_rdata <= 8'hC1;
			14'd5284: ff_rdata <= 8'h67;
			14'd5285: ff_rdata <= 8'hD5;
			14'd5286: ff_rdata <= 8'h7E;
			14'd5287: ff_rdata <= 8'hFE;
			14'd5288: ff_rdata <= 8'h29;
			14'd5289: ff_rdata <= 8'h1E;
			14'd5290: ff_rdata <= 8'h00;
			14'd5291: ff_rdata <= 8'h28;
			14'd5292: ff_rdata <= 8'h06;
			14'd5293: ff_rdata <= 8'hCD;
			14'd5294: ff_rdata <= 8'hDF;
			14'd5295: ff_rdata <= 8'h55;
			14'd5296: ff_rdata <= 8'hCD;
			14'd5297: ff_rdata <= 8'hC1;
			14'd5298: ff_rdata <= 8'h67;
			14'd5299: ff_rdata <= 8'hCD;
			14'd5300: ff_rdata <= 8'hE9;
			14'd5301: ff_rdata <= 8'h55;
			14'd5302: ff_rdata <= 8'h7B;
			14'd5303: ff_rdata <= 8'hB7;
			14'd5304: ff_rdata <= 8'hC2;
			14'd5305: ff_rdata <= 8'h70;
			14'd5306: ff_rdata <= 8'h67;
			14'd5307: ff_rdata <= 8'hD1;
			14'd5308: ff_rdata <= 8'hC1;
			14'd5309: ff_rdata <= 8'h43;
			14'd5310: ff_rdata <= 8'hCD;
			14'd5311: ff_rdata <= 8'hB5;
			14'd5312: ff_rdata <= 8'h6D;
			14'd5313: ff_rdata <= 8'hDA;
			14'd5314: ff_rdata <= 8'h70;
			14'd5315: ff_rdata <= 8'h67;
			14'd5316: ff_rdata <= 8'hC9;
			14'd5317: ff_rdata <= 8'h3E;
			14'd5318: ff_rdata <= 8'h01;
			14'd5319: ff_rdata <= 8'h32;
			14'd5320: ff_rdata <= 8'hA5;
			14'd5321: ff_rdata <= 8'hF6;
			14'd5322: ff_rdata <= 8'hCD;
			14'd5323: ff_rdata <= 8'h9B;
			14'd5324: ff_rdata <= 8'h67;
			14'd5325: ff_rdata <= 8'hC2;
			14'd5326: ff_rdata <= 8'h70;
			14'd5327: ff_rdata <= 8'h67;
			14'd5328: ff_rdata <= 8'h32;
			14'd5329: ff_rdata <= 8'hA5;
			14'd5330: ff_rdata <= 8'hF6;
			14'd5331: ff_rdata <= 8'h3A;
			14'd5332: ff_rdata <= 8'h63;
			14'd5333: ff_rdata <= 8'hF6;
			14'd5334: ff_rdata <= 8'hFE;
			14'd5335: ff_rdata <= 8'h03;
			14'd5336: ff_rdata <= 8'hCA;
			14'd5337: ff_rdata <= 8'h70;
			14'd5338: ff_rdata <= 8'h67;
			14'd5339: ff_rdata <= 8'hEB;
			14'd5340: ff_rdata <= 8'h09;
			14'd5341: ff_rdata <= 8'h2B;
			14'd5342: ff_rdata <= 8'hEB;
			14'd5343: ff_rdata <= 8'h0A;
			14'd5344: ff_rdata <= 8'h37;
			14'd5345: ff_rdata <= 8'h17;
			14'd5346: ff_rdata <= 8'h81;
			14'd5347: ff_rdata <= 8'h4F;
			14'd5348: ff_rdata <= 8'hD0;
			14'd5349: ff_rdata <= 8'h04;
			14'd5350: ff_rdata <= 8'hC9;
			14'd5351: ff_rdata <= 8'h2B;
			14'd5352: ff_rdata <= 8'hC3;
			14'd5353: ff_rdata <= 8'hAF;
			14'd5354: ff_rdata <= 8'h67;
			14'd5355: ff_rdata <= 8'hCD;
			14'd5356: ff_rdata <= 8'hF3;
			14'd5357: ff_rdata <= 8'h54;
			14'd5358: ff_rdata <= 8'hE1;
			14'd5359: ff_rdata <= 8'hCD;
			14'd5360: ff_rdata <= 8'hE9;
			14'd5361: ff_rdata <= 8'h55;
			14'd5362: ff_rdata <= 8'hC9;
			14'd5363: ff_rdata <= 8'h22;
			14'd5364: ff_rdata <= 8'hF8;
			14'd5365: ff_rdata <= 8'hF7;
			14'd5366: ff_rdata <= 8'h21;
			14'd5367: ff_rdata <= 8'h63;
			14'd5368: ff_rdata <= 8'hF6;
			14'd5369: ff_rdata <= 8'h7E;
			14'd5370: ff_rdata <= 8'hFE;
			14'd5371: ff_rdata <= 8'h02;
			14'd5372: ff_rdata <= 8'h28;
			14'd5373: ff_rdata <= 8'h21;
			14'd5374: ff_rdata <= 8'hFE;
			14'd5375: ff_rdata <= 8'h04;
			14'd5376: ff_rdata <= 8'h28;
			14'd5377: ff_rdata <= 8'h0F;
			14'd5378: ff_rdata <= 8'hFE;
			14'd5379: ff_rdata <= 8'h08;
			14'd5380: ff_rdata <= 8'hC2;
			14'd5381: ff_rdata <= 8'h73;
			14'd5382: ff_rdata <= 8'h67;
			14'd5383: ff_rdata <= 8'h36;
			14'd5384: ff_rdata <= 8'h02;
			14'd5385: ff_rdata <= 8'hD5;
			14'd5386: ff_rdata <= 8'hCD;
			14'd5387: ff_rdata <= 8'hA1;
			14'd5388: ff_rdata <= 8'h67;
			14'd5389: ff_rdata <= 8'h0E;
			14'd5390: ff_rdata <= 8'h08;
			14'd5391: ff_rdata <= 8'h18;
			14'd5392: ff_rdata <= 8'h08;
			14'd5393: ff_rdata <= 8'h36;
			14'd5394: ff_rdata <= 8'h02;
			14'd5395: ff_rdata <= 8'hD5;
			14'd5396: ff_rdata <= 8'hCD;
			14'd5397: ff_rdata <= 8'hA1;
			14'd5398: ff_rdata <= 8'h67;
			14'd5399: ff_rdata <= 8'h0E;
			14'd5400: ff_rdata <= 8'h04;
			14'd5401: ff_rdata <= 8'hD1;
			14'd5402: ff_rdata <= 8'h21;
			14'd5403: ff_rdata <= 8'hF6;
			14'd5404: ff_rdata <= 8'hF7;
			14'd5405: ff_rdata <= 8'h18;
			14'd5406: ff_rdata <= 8'h05;
			14'd5407: ff_rdata <= 8'h21;
			14'd5408: ff_rdata <= 8'hF8;
			14'd5409: ff_rdata <= 8'hF7;
			14'd5410: ff_rdata <= 8'h0E;
			14'd5411: ff_rdata <= 8'h02;
			14'd5412: ff_rdata <= 8'h06;
			14'd5413: ff_rdata <= 8'h00;
			14'd5414: ff_rdata <= 8'hED;
			14'd5415: ff_rdata <= 8'hB0;
			14'd5416: ff_rdata <= 8'hC9;
			14'd5417: ff_rdata <= 8'hCD;
			14'd5418: ff_rdata <= 8'h65;
			14'd5419: ff_rdata <= 8'h54;
			14'd5420: ff_rdata <= 8'hE5;
			14'd5421: ff_rdata <= 8'hCD;
			14'd5422: ff_rdata <= 8'h50;
			14'd5423: ff_rdata <= 8'h6B;
			14'd5424: ff_rdata <= 8'hE1;
			14'd5425: ff_rdata <= 8'hDA;
			14'd5426: ff_rdata <= 8'h70;
			14'd5427: ff_rdata <= 8'h67;
			14'd5428: ff_rdata <= 8'hC9;
			14'd5429: ff_rdata <= 8'hCD;
			14'd5430: ff_rdata <= 8'h65;
			14'd5431: ff_rdata <= 8'h54;
			14'd5432: ff_rdata <= 8'hE5;
			14'd5433: ff_rdata <= 8'hCD;
			14'd5434: ff_rdata <= 8'hDA;
			14'd5435: ff_rdata <= 8'h6B;
			14'd5436: ff_rdata <= 8'hE1;
			14'd5437: ff_rdata <= 8'hDA;
			14'd5438: ff_rdata <= 8'h70;
			14'd5439: ff_rdata <= 8'h67;
			14'd5440: ff_rdata <= 8'hC9;
			14'd5441: ff_rdata <= 8'hCD;
			14'd5442: ff_rdata <= 8'hC1;
			14'd5443: ff_rdata <= 8'h52;
			14'd5444: ff_rdata <= 8'h4F;
			14'd5445: ff_rdata <= 8'hCD;
			14'd5446: ff_rdata <= 8'h9F;
			14'd5447: ff_rdata <= 8'h6C;
			14'd5448: ff_rdata <= 8'hDA;
			14'd5449: ff_rdata <= 8'h70;
			14'd5450: ff_rdata <= 8'h67;
			14'd5451: ff_rdata <= 8'hC9;
			14'd5452: ff_rdata <= 8'hC5;
			14'd5453: ff_rdata <= 8'hD5;
			14'd5454: ff_rdata <= 8'hE5;
			14'd5455: ff_rdata <= 8'h06;
			14'd5456: ff_rdata <= 8'h01;
			14'd5457: ff_rdata <= 8'hCD;
			14'd5458: ff_rdata <= 8'h58;
			14'd5459: ff_rdata <= 8'h55;
			14'd5460: ff_rdata <= 8'hE1;
			14'd5461: ff_rdata <= 8'hD1;
			14'd5462: ff_rdata <= 8'hC1;
			14'd5463: ff_rdata <= 8'hC9;
			14'd5464: ff_rdata <= 8'hDB;
			14'd5465: ff_rdata <= 8'hA8;
			14'd5466: ff_rdata <= 8'hCD;
			14'd5467: ff_rdata <= 8'h7A;
			14'd5468: ff_rdata <= 8'h55;
			14'd5469: ff_rdata <= 8'hE6;
			14'd5470: ff_rdata <= 8'h03;
			14'd5471: ff_rdata <= 8'h5F;
			14'd5472: ff_rdata <= 8'h16;
			14'd5473: ff_rdata <= 8'h00;
			14'd5474: ff_rdata <= 8'h21;
			14'd5475: ff_rdata <= 8'hC1;
			14'd5476: ff_rdata <= 8'hFC;
			14'd5477: ff_rdata <= 8'h19;
			14'd5478: ff_rdata <= 8'h7E;
			14'd5479: ff_rdata <= 8'hE6;
			14'd5480: ff_rdata <= 8'h80;
			14'd5481: ff_rdata <= 8'hB3;
			14'd5482: ff_rdata <= 8'hF0;
			14'd5483: ff_rdata <= 8'h5F;
			14'd5484: ff_rdata <= 8'h23;
			14'd5485: ff_rdata <= 8'h23;
			14'd5486: ff_rdata <= 8'h23;
			14'd5487: ff_rdata <= 8'h23;
			14'd5488: ff_rdata <= 8'h7E;
			14'd5489: ff_rdata <= 8'h07;
			14'd5490: ff_rdata <= 8'h07;
			14'd5491: ff_rdata <= 8'hCD;
			14'd5492: ff_rdata <= 8'h7A;
			14'd5493: ff_rdata <= 8'h55;
			14'd5494: ff_rdata <= 8'hE6;
			14'd5495: ff_rdata <= 8'h0C;
			14'd5496: ff_rdata <= 8'hB3;
			14'd5497: ff_rdata <= 8'hC9;
			14'd5498: ff_rdata <= 8'h04;
			14'd5499: ff_rdata <= 8'h05;
			14'd5500: ff_rdata <= 8'hC8;
			14'd5501: ff_rdata <= 8'hC5;
			14'd5502: ff_rdata <= 8'h0F;
			14'd5503: ff_rdata <= 8'h0F;
			14'd5504: ff_rdata <= 8'h10;
			14'd5505: ff_rdata <= 8'hFC;
			14'd5506: ff_rdata <= 8'hC1;
			14'd5507: ff_rdata <= 8'hC9;
			14'd5508: ff_rdata <= 8'hCD;
			14'd5509: ff_rdata <= 8'h61;
			14'd5510: ff_rdata <= 8'h6D;
			14'd5511: ff_rdata <= 8'hDD;
			14'd5512: ff_rdata <= 8'h21;
			14'd5513: ff_rdata <= 8'h27;
			14'd5514: ff_rdata <= 8'hFA;
			14'd5515: ff_rdata <= 8'h01;
			14'd5516: ff_rdata <= 8'h00;
			14'd5517: ff_rdata <= 8'h09;
			14'd5518: ff_rdata <= 8'h79;
			14'd5519: ff_rdata <= 8'hC6;
			14'd5520: ff_rdata <= 8'h10;
			14'd5521: ff_rdata <= 8'hDD;
			14'd5522: ff_rdata <= 8'h77;
			14'd5523: ff_rdata <= 8'h00;
			14'd5524: ff_rdata <= 8'hDD;
			14'd5525: ff_rdata <= 8'h36;
			14'd5526: ff_rdata <= 8'h01;
			14'd5527: ff_rdata <= 8'h04;
			14'd5528: ff_rdata <= 8'hDD;
			14'd5529: ff_rdata <= 8'h36;
			14'd5530: ff_rdata <= 8'h02;
			14'd5531: ff_rdata <= 8'h00;
			14'd5532: ff_rdata <= 8'hDD;
			14'd5533: ff_rdata <= 8'h36;
			14'd5534: ff_rdata <= 8'h03;
			14'd5535: ff_rdata <= 8'h00;
			14'd5536: ff_rdata <= 8'hDD;
			14'd5537: ff_rdata <= 8'h36;
			14'd5538: ff_rdata <= 8'h04;
			14'd5539: ff_rdata <= 8'h00;
			14'd5540: ff_rdata <= 8'hDD;
			14'd5541: ff_rdata <= 8'h36;
			14'd5542: ff_rdata <= 8'h05;
			14'd5543: ff_rdata <= 8'h00;
			14'd5544: ff_rdata <= 8'hDD;
			14'd5545: ff_rdata <= 8'h36;
			14'd5546: ff_rdata <= 8'h06;
			14'd5547: ff_rdata <= 8'h00;
			14'd5548: ff_rdata <= 8'h11;
			14'd5549: ff_rdata <= 8'h10;
			14'd5550: ff_rdata <= 8'h00;
			14'd5551: ff_rdata <= 8'hDD;
			14'd5552: ff_rdata <= 8'h19;
			14'd5553: ff_rdata <= 8'h0C;
			14'd5554: ff_rdata <= 8'h10;
			14'd5555: ff_rdata <= 8'hDA;
			14'd5556: ff_rdata <= 8'h3A;
			14'd5557: ff_rdata <= 8'h8E;
			14'd5558: ff_rdata <= 8'hF9;
			14'd5559: ff_rdata <= 8'hE6;
			14'd5560: ff_rdata <= 8'h01;
			14'd5561: ff_rdata <= 8'hC4;
			14'd5562: ff_rdata <= 8'h86;
			14'd5563: ff_rdata <= 8'h6D;
			14'd5564: ff_rdata <= 8'h0E;
			14'd5565: ff_rdata <= 8'h09;
			14'd5566: ff_rdata <= 8'hCD;
			14'd5567: ff_rdata <= 8'h9F;
			14'd5568: ff_rdata <= 8'h6C;
			14'd5569: ff_rdata <= 8'hDD;
			14'd5570: ff_rdata <= 8'h21;
			14'd5571: ff_rdata <= 8'h27;
			14'd5572: ff_rdata <= 8'hFA;
			14'd5573: ff_rdata <= 8'h3A;
			14'd5574: ff_rdata <= 8'h8E;
			14'd5575: ff_rdata <= 8'hF9;
			14'd5576: ff_rdata <= 8'hE6;
			14'd5577: ff_rdata <= 8'h01;
			14'd5578: ff_rdata <= 8'h06;
			14'd5579: ff_rdata <= 8'h09;
			14'd5580: ff_rdata <= 8'h28;
			14'd5581: ff_rdata <= 8'h02;
			14'd5582: ff_rdata <= 8'h06;
			14'd5583: ff_rdata <= 8'h06;
			14'd5584: ff_rdata <= 8'hC5;
			14'd5585: ff_rdata <= 8'h0E;
			14'd5586: ff_rdata <= 8'h00;
			14'd5587: ff_rdata <= 8'hCD;
			14'd5588: ff_rdata <= 8'hE1;
			14'd5589: ff_rdata <= 8'h68;
			14'd5590: ff_rdata <= 8'hC1;
			14'd5591: ff_rdata <= 8'h11;
			14'd5592: ff_rdata <= 8'h10;
			14'd5593: ff_rdata <= 8'h00;
			14'd5594: ff_rdata <= 8'hDD;
			14'd5595: ff_rdata <= 8'h19;
			14'd5596: ff_rdata <= 8'h10;
			14'd5597: ff_rdata <= 8'hF2;
			14'd5598: ff_rdata <= 8'hC9;
			14'd5599: ff_rdata <= 8'hCD;
			14'd5600: ff_rdata <= 8'hA7;
			14'd5601: ff_rdata <= 8'h67;
			14'd5602: ff_rdata <= 8'h2C;
			14'd5603: ff_rdata <= 8'hC9;
			14'd5604: ff_rdata <= 8'hCD;
			14'd5605: ff_rdata <= 8'hA7;
			14'd5606: ff_rdata <= 8'h67;
			14'd5607: ff_rdata <= 8'h28;
			14'd5608: ff_rdata <= 8'hC9;
			14'd5609: ff_rdata <= 8'hCD;
			14'd5610: ff_rdata <= 8'hA7;
			14'd5611: ff_rdata <= 8'h67;
			14'd5612: ff_rdata <= 8'h29;
			14'd5613: ff_rdata <= 8'hC9;
			14'd5614: ff_rdata <= 8'hCD;
			14'd5615: ff_rdata <= 8'hA7;
			14'd5616: ff_rdata <= 8'h67;
			14'd5617: ff_rdata <= 8'h28;
			14'd5618: ff_rdata <= 8'h11;
			14'd5619: ff_rdata <= 8'h5E;
			14'd5620: ff_rdata <= 8'hF5;
			14'd5621: ff_rdata <= 8'h06;
			14'd5622: ff_rdata <= 8'h09;
			14'd5623: ff_rdata <= 8'h7E;
			14'd5624: ff_rdata <= 8'hFE;
			14'd5625: ff_rdata <= 8'h2C;
			14'd5626: ff_rdata <= 8'h28;
			14'd5627: ff_rdata <= 8'h1F;
			14'd5628: ff_rdata <= 8'hC5;
			14'd5629: ff_rdata <= 8'h3E;
			14'd5630: ff_rdata <= 8'h09;
			14'd5631: ff_rdata <= 8'h90;
			14'd5632: ff_rdata <= 8'h12;
			14'd5633: ff_rdata <= 8'h13;
			14'd5634: ff_rdata <= 8'hD5;
			14'd5635: ff_rdata <= 8'h7E;
			14'd5636: ff_rdata <= 8'hCD;
			14'd5637: ff_rdata <= 8'hC5;
			14'd5638: ff_rdata <= 8'h56;
			14'd5639: ff_rdata <= 8'h3E;
			14'd5640: ff_rdata <= 8'h00;
			14'd5641: ff_rdata <= 8'h38;
			14'd5642: ff_rdata <= 8'h01;
			14'd5643: ff_rdata <= 8'h2F;
			14'd5644: ff_rdata <= 8'hE3;
			14'd5645: ff_rdata <= 8'h77;
			14'd5646: ff_rdata <= 8'h23;
			14'd5647: ff_rdata <= 8'h73;
			14'd5648: ff_rdata <= 8'h23;
			14'd5649: ff_rdata <= 8'h72;
			14'd5650: ff_rdata <= 8'h23;
			14'd5651: ff_rdata <= 8'hE3;
			14'd5652: ff_rdata <= 8'hD1;
			14'd5653: ff_rdata <= 8'hC1;
			14'd5654: ff_rdata <= 8'h7E;
			14'd5655: ff_rdata <= 8'hFE;
			14'd5656: ff_rdata <= 8'h29;
			14'd5657: ff_rdata <= 8'h28;
			14'd5658: ff_rdata <= 8'h06;
			14'd5659: ff_rdata <= 8'hCD;
			14'd5660: ff_rdata <= 8'hA7;
			14'd5661: ff_rdata <= 8'h67;
			14'd5662: ff_rdata <= 8'h2C;
			14'd5663: ff_rdata <= 8'h10;
			14'd5664: ff_rdata <= 8'hD6;
			14'd5665: ff_rdata <= 8'hCD;
			14'd5666: ff_rdata <= 8'hA7;
			14'd5667: ff_rdata <= 8'h67;
			14'd5668: ff_rdata <= 8'h29;
			14'd5669: ff_rdata <= 8'hC2;
			14'd5670: ff_rdata <= 8'h6D;
			14'd5671: ff_rdata <= 8'h67;
			14'd5672: ff_rdata <= 8'h3E;
			14'd5673: ff_rdata <= 8'hFF;
			14'd5674: ff_rdata <= 8'h12;
			14'd5675: ff_rdata <= 8'hCD;
			14'd5676: ff_rdata <= 8'h32;
			14'd5677: ff_rdata <= 8'h56;
			14'd5678: ff_rdata <= 8'hDA;
			14'd5679: ff_rdata <= 8'h70;
			14'd5680: ff_rdata <= 8'h67;
			14'd5681: ff_rdata <= 8'hC9;
			14'd5682: ff_rdata <= 8'hE5;
			14'd5683: ff_rdata <= 8'h21;
			14'd5684: ff_rdata <= 8'h5E;
			14'd5685: ff_rdata <= 8'hF5;
			14'd5686: ff_rdata <= 8'h7E;
			14'd5687: ff_rdata <= 8'hFE;
			14'd5688: ff_rdata <= 8'hFF;
			14'd5689: ff_rdata <= 8'h28;
			14'd5690: ff_rdata <= 8'h27;
			14'd5691: ff_rdata <= 8'h23;
			14'd5692: ff_rdata <= 8'hCD;
			14'd5693: ff_rdata <= 8'h6D;
			14'd5694: ff_rdata <= 8'h56;
			14'd5695: ff_rdata <= 8'h7E;
			14'd5696: ff_rdata <= 8'h23;
			14'd5697: ff_rdata <= 8'hB7;
			14'd5698: ff_rdata <= 8'h28;
			14'd5699: ff_rdata <= 8'h0C;
			14'd5700: ff_rdata <= 8'h4E;
			14'd5701: ff_rdata <= 8'h23;
			14'd5702: ff_rdata <= 8'h46;
			14'd5703: ff_rdata <= 8'hE5;
			14'd5704: ff_rdata <= 8'hCD;
			14'd5705: ff_rdata <= 8'hDA;
			14'd5706: ff_rdata <= 8'h68;
			14'd5707: ff_rdata <= 8'hCD;
			14'd5708: ff_rdata <= 8'h65;
			14'd5709: ff_rdata <= 8'h56;
			14'd5710: ff_rdata <= 8'h18;
			14'd5711: ff_rdata <= 8'h0E;
			14'd5712: ff_rdata <= 8'h4E;
			14'd5713: ff_rdata <= 8'h79;
			14'd5714: ff_rdata <= 8'hFE;
			14'd5715: ff_rdata <= 8'h40;
			14'd5716: ff_rdata <= 8'h3F;
			14'd5717: ff_rdata <= 8'hD8;
			14'd5718: ff_rdata <= 8'h23;
			14'd5719: ff_rdata <= 8'hE5;
			14'd5720: ff_rdata <= 8'hCD;
			14'd5721: ff_rdata <= 8'hE1;
			14'd5722: ff_rdata <= 8'h68;
			14'd5723: ff_rdata <= 8'hCD;
			14'd5724: ff_rdata <= 8'h65;
			14'd5725: ff_rdata <= 8'h56;
			14'd5726: ff_rdata <= 8'hE1;
			14'd5727: ff_rdata <= 8'h23;
			14'd5728: ff_rdata <= 8'h18;
			14'd5729: ff_rdata <= 8'hD4;
			14'd5730: ff_rdata <= 8'hE1;
			14'd5731: ff_rdata <= 8'hB7;
			14'd5732: ff_rdata <= 8'hC9;
			14'd5733: ff_rdata <= 8'hC5;
			14'd5734: ff_rdata <= 8'h01;
			14'd5735: ff_rdata <= 8'h10;
			14'd5736: ff_rdata <= 8'h00;
			14'd5737: ff_rdata <= 8'hDD;
			14'd5738: ff_rdata <= 8'h09;
			14'd5739: ff_rdata <= 8'hC1;
			14'd5740: ff_rdata <= 8'hC9;
			14'd5741: ff_rdata <= 8'hDD;
			14'd5742: ff_rdata <= 8'h21;
			14'd5743: ff_rdata <= 8'h27;
			14'd5744: ff_rdata <= 8'hFA;
			14'd5745: ff_rdata <= 8'hB7;
			14'd5746: ff_rdata <= 8'hC8;
			14'd5747: ff_rdata <= 8'hC5;
			14'd5748: ff_rdata <= 8'h01;
			14'd5749: ff_rdata <= 8'h10;
			14'd5750: ff_rdata <= 8'h00;
			14'd5751: ff_rdata <= 8'hDD;
			14'd5752: ff_rdata <= 8'h09;
			14'd5753: ff_rdata <= 8'h3D;
			14'd5754: ff_rdata <= 8'h20;
			14'd5755: ff_rdata <= 8'hFB;
			14'd5756: ff_rdata <= 8'hC1;
			14'd5757: ff_rdata <= 8'hC9;
			14'd5758: ff_rdata <= 8'hCD;
			14'd5759: ff_rdata <= 8'hA7;
			14'd5760: ff_rdata <= 8'h67;
			14'd5761: ff_rdata <= 8'h28;
			14'd5762: ff_rdata <= 8'hCD;
			14'd5763: ff_rdata <= 8'hC5;
			14'd5764: ff_rdata <= 8'h56;
			14'd5765: ff_rdata <= 8'h3F;
			14'd5766: ff_rdata <= 8'h9F;
			14'd5767: ff_rdata <= 8'h32;
			14'd5768: ff_rdata <= 8'h5E;
			14'd5769: ff_rdata <= 8'hF5;
			14'd5770: ff_rdata <= 8'hED;
			14'd5771: ff_rdata <= 8'h53;
			14'd5772: ff_rdata <= 8'h5F;
			14'd5773: ff_rdata <= 8'hF5;
			14'd5774: ff_rdata <= 8'hED;
			14'd5775: ff_rdata <= 8'h43;
			14'd5776: ff_rdata <= 8'h61;
			14'd5777: ff_rdata <= 8'hF5;
			14'd5778: ff_rdata <= 8'hCD;
			14'd5779: ff_rdata <= 8'hA7;
			14'd5780: ff_rdata <= 8'h67;
			14'd5781: ff_rdata <= 8'h2C;
			14'd5782: ff_rdata <= 8'hCD;
			14'd5783: ff_rdata <= 8'hC5;
			14'd5784: ff_rdata <= 8'h56;
			14'd5785: ff_rdata <= 8'h3F;
			14'd5786: ff_rdata <= 8'h9F;
			14'd5787: ff_rdata <= 8'h32;
			14'd5788: ff_rdata <= 8'h63;
			14'd5789: ff_rdata <= 8'hF5;
			14'd5790: ff_rdata <= 8'hED;
			14'd5791: ff_rdata <= 8'h53;
			14'd5792: ff_rdata <= 8'h64;
			14'd5793: ff_rdata <= 8'hF5;
			14'd5794: ff_rdata <= 8'hED;
			14'd5795: ff_rdata <= 8'h43;
			14'd5796: ff_rdata <= 8'h66;
			14'd5797: ff_rdata <= 8'hF5;
			14'd5798: ff_rdata <= 8'h20;
			14'd5799: ff_rdata <= 8'h05;
			14'd5800: ff_rdata <= 8'h7B;
			14'd5801: ff_rdata <= 8'hFE;
			14'd5802: ff_rdata <= 8'h20;
			14'd5803: ff_rdata <= 8'h38;
			14'd5804: ff_rdata <= 8'h31;
			14'd5805: ff_rdata <= 8'hCD;
			14'd5806: ff_rdata <= 8'hA7;
			14'd5807: ff_rdata <= 8'h67;
			14'd5808: ff_rdata <= 8'h29;
			14'd5809: ff_rdata <= 8'hC2;
			14'd5810: ff_rdata <= 8'h6D;
			14'd5811: ff_rdata <= 8'h67;
			14'd5812: ff_rdata <= 8'hE5;
			14'd5813: ff_rdata <= 8'h21;
			14'd5814: ff_rdata <= 8'h5E;
			14'd5815: ff_rdata <= 8'hF5;
			14'd5816: ff_rdata <= 8'h3A;
			14'd5817: ff_rdata <= 8'h63;
			14'd5818: ff_rdata <= 8'hF5;
			14'd5819: ff_rdata <= 8'hA6;
			14'd5820: ff_rdata <= 8'h20;
			14'd5821: ff_rdata <= 8'h20;
			14'd5822: ff_rdata <= 8'hCD;
			14'd5823: ff_rdata <= 8'hF9;
			14'd5824: ff_rdata <= 8'h56;
			14'd5825: ff_rdata <= 8'h38;
			14'd5826: ff_rdata <= 8'h1B;
			14'd5827: ff_rdata <= 8'hE1;
			14'd5828: ff_rdata <= 8'hC9;
			14'd5829: ff_rdata <= 8'hFE;
			14'd5830: ff_rdata <= 8'h40;
			14'd5831: ff_rdata <= 8'h28;
			14'd5832: ff_rdata <= 8'h0C;
			14'd5833: ff_rdata <= 8'hFE;
			14'd5834: ff_rdata <= 8'hF3;
			14'd5835: ff_rdata <= 8'h20;
			14'd5836: ff_rdata <= 8'h14;
			14'd5837: ff_rdata <= 8'hCD;
			14'd5838: ff_rdata <= 8'hAF;
			14'd5839: ff_rdata <= 8'h67;
			14'd5840: ff_rdata <= 8'h11;
			14'd5841: ff_rdata <= 8'hFF;
			14'd5842: ff_rdata <= 8'h00;
			14'd5843: ff_rdata <= 8'h37;
			14'd5844: ff_rdata <= 8'hC9;
			14'd5845: ff_rdata <= 8'hCD;
			14'd5846: ff_rdata <= 8'hAF;
			14'd5847: ff_rdata <= 8'h67;
			14'd5848: ff_rdata <= 8'hCD;
			14'd5849: ff_rdata <= 8'hC1;
			14'd5850: ff_rdata <= 8'h67;
			14'd5851: ff_rdata <= 8'hFE;
			14'd5852: ff_rdata <= 8'h40;
			14'd5853: ff_rdata <= 8'hD8;
			14'd5854: ff_rdata <= 8'hC3;
			14'd5855: ff_rdata <= 8'h70;
			14'd5856: ff_rdata <= 8'h67;
			14'd5857: ff_rdata <= 8'hCD;
			14'd5858: ff_rdata <= 8'hEF;
			14'd5859: ff_rdata <= 8'h56;
			14'd5860: ff_rdata <= 8'h7B;
			14'd5861: ff_rdata <= 8'hE6;
			14'd5862: ff_rdata <= 8'hE0;
			14'd5863: ff_rdata <= 8'hB2;
			14'd5864: ff_rdata <= 8'h28;
			14'd5865: ff_rdata <= 8'hF4;
			14'd5866: ff_rdata <= 8'hD5;
			14'd5867: ff_rdata <= 8'h59;
			14'd5868: ff_rdata <= 8'h50;
			14'd5869: ff_rdata <= 8'hC1;
			14'd5870: ff_rdata <= 8'hC9;
			14'd5871: ff_rdata <= 8'hCD;
			14'd5872: ff_rdata <= 8'hC5;
			14'd5873: ff_rdata <= 8'h54;
			14'd5874: ff_rdata <= 8'hEB;
			14'd5875: ff_rdata <= 8'hB7;
			14'd5876: ff_rdata <= 8'hED;
			14'd5877: ff_rdata <= 8'h42;
			14'd5878: ff_rdata <= 8'h23;
			14'd5879: ff_rdata <= 8'hEB;
			14'd5880: ff_rdata <= 8'hC9;
			14'd5881: ff_rdata <= 8'h3A;
			14'd5882: ff_rdata <= 8'h63;
			14'd5883: ff_rdata <= 8'hF5;
			14'd5884: ff_rdata <= 8'h2A;
			14'd5885: ff_rdata <= 8'h64;
			14'd5886: ff_rdata <= 8'hF5;
			14'd5887: ff_rdata <= 8'hB7;
			14'd5888: ff_rdata <= 8'h20;
			14'd5889: ff_rdata <= 8'h0B;
			14'd5890: ff_rdata <= 8'h7D;
			14'd5891: ff_rdata <= 8'h3C;
			14'd5892: ff_rdata <= 8'h37;
			14'd5893: ff_rdata <= 8'hC8;
			14'd5894: ff_rdata <= 8'hFE;
			14'd5895: ff_rdata <= 8'h40;
			14'd5896: ff_rdata <= 8'h37;
			14'd5897: ff_rdata <= 8'hC0;
			14'd5898: ff_rdata <= 8'h21;
			14'd5899: ff_rdata <= 8'hF9;
			14'd5900: ff_rdata <= 8'hF9;
			14'd5901: ff_rdata <= 8'hE5;
			14'd5902: ff_rdata <= 8'h3A;
			14'd5903: ff_rdata <= 8'h5E;
			14'd5904: ff_rdata <= 8'hF5;
			14'd5905: ff_rdata <= 8'h2A;
			14'd5906: ff_rdata <= 8'h5F;
			14'd5907: ff_rdata <= 8'hF5;
			14'd5908: ff_rdata <= 8'hB7;
			14'd5909: ff_rdata <= 8'h20;
			14'd5910: ff_rdata <= 8'h0E;
			14'd5911: ff_rdata <= 8'h7D;
			14'd5912: ff_rdata <= 8'hFE;
			14'd5913: ff_rdata <= 8'hFF;
			14'd5914: ff_rdata <= 8'h28;
			14'd5915: ff_rdata <= 8'h13;
			14'd5916: ff_rdata <= 8'h4F;
			14'd5917: ff_rdata <= 8'hCD;
			14'd5918: ff_rdata <= 8'h0F;
			14'd5919: ff_rdata <= 8'h69;
			14'd5920: ff_rdata <= 8'h28;
			14'd5921: ff_rdata <= 8'h0D;
			14'd5922: ff_rdata <= 8'hCD;
			14'd5923: ff_rdata <= 8'h32;
			14'd5924: ff_rdata <= 8'h57;
			14'd5925: ff_rdata <= 8'hD1;
			14'd5926: ff_rdata <= 8'h01;
			14'd5927: ff_rdata <= 8'h20;
			14'd5928: ff_rdata <= 8'h00;
			14'd5929: ff_rdata <= 8'hF3;
			14'd5930: ff_rdata <= 8'hED;
			14'd5931: ff_rdata <= 8'hB0;
			14'd5932: ff_rdata <= 8'hB7;
			14'd5933: ff_rdata <= 8'hFB;
			14'd5934: ff_rdata <= 8'hC9;
			14'd5935: ff_rdata <= 8'hE1;
			14'd5936: ff_rdata <= 8'h37;
			14'd5937: ff_rdata <= 8'hC9;
			14'd5938: ff_rdata <= 8'h7D;
			14'd5939: ff_rdata <= 8'hFE;
			14'd5940: ff_rdata <= 8'h3F;
			14'd5941: ff_rdata <= 8'h21;
			14'd5942: ff_rdata <= 8'hF9;
			14'd5943: ff_rdata <= 8'hF9;
			14'd5944: ff_rdata <= 8'hC8;
			14'd5945: ff_rdata <= 8'h6F;
			14'd5946: ff_rdata <= 8'h26;
			14'd5947: ff_rdata <= 8'h00;
			14'd5948: ff_rdata <= 8'h29;
			14'd5949: ff_rdata <= 8'h29;
			14'd5950: ff_rdata <= 8'h29;
			14'd5951: ff_rdata <= 8'h29;
			14'd5952: ff_rdata <= 8'h29;
			14'd5953: ff_rdata <= 8'h11;
			14'd5954: ff_rdata <= 8'h0C;
			14'd5955: ff_rdata <= 8'h6E;
			14'd5956: ff_rdata <= 8'h19;
			14'd5957: ff_rdata <= 8'hC9;
			14'd5958: ff_rdata <= 8'hCD;
			14'd5959: ff_rdata <= 8'hB4;
			14'd5960: ff_rdata <= 8'h52;
			14'd5961: ff_rdata <= 8'h3A;
			14'd5962: ff_rdata <= 8'h91;
			14'd5963: ff_rdata <= 8'hF9;
			14'd5964: ff_rdata <= 8'hBB;
			14'd5965: ff_rdata <= 8'hDA;
			14'd5966: ff_rdata <= 8'h70;
			14'd5967: ff_rdata <= 8'h67;
			14'd5968: ff_rdata <= 8'h7B;
			14'd5969: ff_rdata <= 8'hE5;
			14'd5970: ff_rdata <= 8'hCD;
			14'd5971: ff_rdata <= 8'h60;
			14'd5972: ff_rdata <= 8'h57;
			14'd5973: ff_rdata <= 8'hE3;
			14'd5974: ff_rdata <= 8'hCD;
			14'd5975: ff_rdata <= 8'hDF;
			14'd5976: ff_rdata <= 8'h55;
			14'd5977: ff_rdata <= 8'hCD;
			14'd5978: ff_rdata <= 8'h9B;
			14'd5979: ff_rdata <= 8'h67;
			14'd5980: ff_rdata <= 8'hE3;
			14'd5981: ff_rdata <= 8'hC3;
			14'd5982: ff_rdata <= 8'hEB;
			14'd5983: ff_rdata <= 8'h54;
			14'd5984: ff_rdata <= 8'h2A;
			14'd5985: ff_rdata <= 8'h95;
			14'd5986: ff_rdata <= 8'hF9;
			14'd5987: ff_rdata <= 8'hB7;
			14'd5988: ff_rdata <= 8'h20;
			14'd5989: ff_rdata <= 8'h0B;
			14'd5990: ff_rdata <= 8'h7C;
			14'd5991: ff_rdata <= 8'hE6;
			14'd5992: ff_rdata <= 8'h1F;
			14'd5993: ff_rdata <= 8'hB5;
			14'd5994: ff_rdata <= 8'h28;
			14'd5995: ff_rdata <= 8'h02;
			14'd5996: ff_rdata <= 8'h3E;
			14'd5997: ff_rdata <= 8'hFF;
			14'd5998: ff_rdata <= 8'h6F;
			14'd5999: ff_rdata <= 8'h67;
			14'd6000: ff_rdata <= 8'hC9;
			14'd6001: ff_rdata <= 8'hCB;
			14'd6002: ff_rdata <= 8'h3C;
			14'd6003: ff_rdata <= 8'hCB;
			14'd6004: ff_rdata <= 8'h1D;
			14'd6005: ff_rdata <= 8'h3D;
			14'd6006: ff_rdata <= 8'h20;
			14'd6007: ff_rdata <= 8'hF9;
			14'd6008: ff_rdata <= 8'h9F;
			14'd6009: ff_rdata <= 8'h18;
			14'd6010: ff_rdata <= 8'hF3;
			14'd6011: ff_rdata <= 8'h3A;
			14'd6012: ff_rdata <= 8'h7C;
			14'd6013: ff_rdata <= 8'hF9;
			14'd6014: ff_rdata <= 8'hF5;
			14'd6015: ff_rdata <= 8'hC5;
			14'd6016: ff_rdata <= 8'hD5;
			14'd6017: ff_rdata <= 8'hE5;
			14'd6018: ff_rdata <= 8'h3A;
			14'd6019: ff_rdata <= 8'hC1;
			14'd6020: ff_rdata <= 8'hFC;
			14'd6021: ff_rdata <= 8'h26;
			14'd6022: ff_rdata <= 8'h40;
			14'd6023: ff_rdata <= 8'hCD;
			14'd6024: ff_rdata <= 8'h24;
			14'd6025: ff_rdata <= 8'h00;
			14'd6026: ff_rdata <= 8'hE1;
			14'd6027: ff_rdata <= 8'hD1;
			14'd6028: ff_rdata <= 8'hC1;
			14'd6029: ff_rdata <= 8'hCD;
			14'd6030: ff_rdata <= 8'h8A;
			14'd6031: ff_rdata <= 8'h2F;
			14'd6032: ff_rdata <= 8'hF1;
			14'd6033: ff_rdata <= 8'hF5;
			14'd6034: ff_rdata <= 8'hC5;
			14'd6035: ff_rdata <= 8'hD5;
			14'd6036: ff_rdata <= 8'hE5;
			14'd6037: ff_rdata <= 8'h26;
			14'd6038: ff_rdata <= 8'h40;
			14'd6039: ff_rdata <= 8'hCD;
			14'd6040: ff_rdata <= 8'h24;
			14'd6041: ff_rdata <= 8'h00;
			14'd6042: ff_rdata <= 8'hE1;
			14'd6043: ff_rdata <= 8'hD1;
			14'd6044: ff_rdata <= 8'hC1;
			14'd6045: ff_rdata <= 8'hF1;
			14'd6046: ff_rdata <= 8'hFB;
			14'd6047: ff_rdata <= 8'hC9;
			14'd6048: ff_rdata <= 8'h20;
			14'd6049: ff_rdata <= 8'hCD;
			14'd6050: ff_rdata <= 8'h0F;
			14'd6051: ff_rdata <= 8'h51;
			14'd6052: ff_rdata <= 8'hCD;
			14'd6053: ff_rdata <= 8'hD9;
			14'd6054: ff_rdata <= 8'h57;
			14'd6055: ff_rdata <= 8'hE5;
			14'd6056: ff_rdata <= 8'h3A;
			14'd6057: ff_rdata <= 8'h7C;
			14'd6058: ff_rdata <= 8'hF9;
			14'd6059: ff_rdata <= 8'hF3;
			14'd6060: ff_rdata <= 8'h87;
			14'd6061: ff_rdata <= 8'h21;
			14'd6062: ff_rdata <= 8'h08;
			14'd6063: ff_rdata <= 8'h00;
			14'd6064: ff_rdata <= 8'h30;
			14'd6065: ff_rdata <= 8'h02;
			14'd6066: ff_rdata <= 8'h2E;
			14'd6067: ff_rdata <= 8'h10;
			14'd6068: ff_rdata <= 8'h39;
			14'd6069: ff_rdata <= 8'hE5;
			14'd6070: ff_rdata <= 8'h5E;
			14'd6071: ff_rdata <= 8'h23;
			14'd6072: ff_rdata <= 8'h56;
			14'd6073: ff_rdata <= 8'h21;
			14'd6074: ff_rdata <= 8'hE8;
			14'd6075: ff_rdata <= 8'h73;
			14'd6076: ff_rdata <= 8'hB7;
			14'd6077: ff_rdata <= 8'hED;
			14'd6078: ff_rdata <= 8'h52;
			14'd6079: ff_rdata <= 8'hC2;
			14'd6080: ff_rdata <= 8'h64;
			14'd6081: ff_rdata <= 8'h67;
			14'd6082: ff_rdata <= 8'hE1;
			14'd6083: ff_rdata <= 8'h2B;
			14'd6084: ff_rdata <= 8'h54;
			14'd6085: ff_rdata <= 8'h5D;
			14'd6086: ff_rdata <= 8'h13;
			14'd6087: ff_rdata <= 8'h13;
			14'd6088: ff_rdata <= 8'h3A;
			14'd6089: ff_rdata <= 8'h7C;
			14'd6090: ff_rdata <= 8'hF9;
			14'd6091: ff_rdata <= 8'h87;
			14'd6092: ff_rdata <= 8'h01;
			14'd6093: ff_rdata <= 8'h08;
			14'd6094: ff_rdata <= 8'h00;
			14'd6095: ff_rdata <= 8'h30;
			14'd6096: ff_rdata <= 8'h02;
			14'd6097: ff_rdata <= 8'h0E;
			14'd6098: ff_rdata <= 8'h10;
			14'd6099: ff_rdata <= 8'hED;
			14'd6100: ff_rdata <= 8'hB8;
			14'd6101: ff_rdata <= 8'hFB;
			14'd6102: ff_rdata <= 8'hE1;
			14'd6103: ff_rdata <= 8'hE1;
			14'd6104: ff_rdata <= 8'hC9;
			14'd6105: ff_rdata <= 8'hFE;
			14'd6106: ff_rdata <= 8'h23;
			14'd6107: ff_rdata <= 8'h20;
			14'd6108: ff_rdata <= 8'h1B;
			14'd6109: ff_rdata <= 8'hCD;
			14'd6110: ff_rdata <= 8'hAF;
			14'd6111: ff_rdata <= 8'h67;
			14'd6112: ff_rdata <= 8'hCD;
			14'd6113: ff_rdata <= 8'hC1;
			14'd6114: ff_rdata <= 8'h67;
			14'd6115: ff_rdata <= 8'hF5;
			14'd6116: ff_rdata <= 8'hCD;
			14'd6117: ff_rdata <= 8'hDF;
			14'd6118: ff_rdata <= 8'h55;
			14'd6119: ff_rdata <= 8'hF1;
			14'd6120: ff_rdata <= 8'hB7;
			14'd6121: ff_rdata <= 8'h28;
			14'd6122: ff_rdata <= 8'h0D;
			14'd6123: ff_rdata <= 8'h3D;
			14'd6124: ff_rdata <= 8'h28;
			14'd6125: ff_rdata <= 8'h04;
			14'd6126: ff_rdata <= 8'hD6;
			14'd6127: ff_rdata <= 8'h03;
			14'd6128: ff_rdata <= 8'h38;
			14'd6129: ff_rdata <= 8'h39;
			14'd6130: ff_rdata <= 8'hC3;
			14'd6131: ff_rdata <= 8'h70;
			14'd6132: ff_rdata <= 8'h67;
			14'd6133: ff_rdata <= 8'h3C;
			14'd6134: ff_rdata <= 8'h18;
			14'd6135: ff_rdata <= 8'h34;
			14'd6136: ff_rdata <= 8'hAF;
			14'd6137: ff_rdata <= 8'h32;
			14'd6138: ff_rdata <= 8'h7F;
			14'd6139: ff_rdata <= 8'hF9;
			14'd6140: ff_rdata <= 8'hE5;
			14'd6141: ff_rdata <= 8'h3A;
			14'd6142: ff_rdata <= 8'h92;
			14'd6143: ff_rdata <= 8'hF9;
			14'd6144: ff_rdata <= 8'hB7;
			14'd6145: ff_rdata <= 8'h28;
			14'd6146: ff_rdata <= 8'h1E;
			14'd6147: ff_rdata <= 8'h47;
			14'd6148: ff_rdata <= 8'hC5;
			14'd6149: ff_rdata <= 8'h78;
			14'd6150: ff_rdata <= 8'h3D;
			14'd6151: ff_rdata <= 8'hCD;
			14'd6152: ff_rdata <= 8'hE0;
			14'd6153: ff_rdata <= 8'h67;
			14'd6154: ff_rdata <= 8'h11;
			14'd6155: ff_rdata <= 8'hA0;
			14'd6156: ff_rdata <= 8'h57;
			14'd6157: ff_rdata <= 8'h36;
			14'd6158: ff_rdata <= 8'h01;
			14'd6159: ff_rdata <= 8'h23;
			14'd6160: ff_rdata <= 8'h73;
			14'd6161: ff_rdata <= 8'h23;
			14'd6162: ff_rdata <= 8'h72;
			14'd6163: ff_rdata <= 8'h23;
			14'd6164: ff_rdata <= 8'h54;
			14'd6165: ff_rdata <= 8'h5D;
			14'd6166: ff_rdata <= 8'h01;
			14'd6167: ff_rdata <= 8'h1C;
			14'd6168: ff_rdata <= 8'h00;
			14'd6169: ff_rdata <= 8'h09;
			14'd6170: ff_rdata <= 8'hEB;
			14'd6171: ff_rdata <= 8'h73;
			14'd6172: ff_rdata <= 8'h23;
			14'd6173: ff_rdata <= 8'h72;
			14'd6174: ff_rdata <= 8'hC1;
			14'd6175: ff_rdata <= 8'h10;
			14'd6176: ff_rdata <= 8'hE3;
			14'd6177: ff_rdata <= 8'hE1;
			14'd6178: ff_rdata <= 8'hAF;
			14'd6179: ff_rdata <= 8'h32;
			14'd6180: ff_rdata <= 8'h35;
			14'd6181: ff_rdata <= 8'hFB;
			14'd6182: ff_rdata <= 8'h3A;
			14'd6183: ff_rdata <= 8'h92;
			14'd6184: ff_rdata <= 8'hF9;
			14'd6185: ff_rdata <= 8'h18;
			14'd6186: ff_rdata <= 8'h08;
			14'd6187: ff_rdata <= 8'hAF;
			14'd6188: ff_rdata <= 8'h32;
			14'd6189: ff_rdata <= 8'h7F;
			14'd6190: ff_rdata <= 8'hF9;
			14'd6191: ff_rdata <= 8'hAF;
			14'd6192: ff_rdata <= 8'h32;
			14'd6193: ff_rdata <= 8'h35;
			14'd6194: ff_rdata <= 8'hFB;
			14'd6195: ff_rdata <= 8'hE5;
			14'd6196: ff_rdata <= 8'h21;
			14'd6197: ff_rdata <= 8'hF6;
			14'd6198: ff_rdata <= 8'hFF;
			14'd6199: ff_rdata <= 8'h39;
			14'd6200: ff_rdata <= 8'h22;
			14'd6201: ff_rdata <= 8'h36;
			14'd6202: ff_rdata <= 8'hFB;
			14'd6203: ff_rdata <= 8'hE1;
			14'd6204: ff_rdata <= 8'hF5;
			14'd6205: ff_rdata <= 8'hE5;
			14'd6206: ff_rdata <= 8'h21;
			14'd6207: ff_rdata <= 8'h7B;
			14'd6208: ff_rdata <= 8'h57;
			14'd6209: ff_rdata <= 8'h11;
			14'd6210: ff_rdata <= 8'hDE;
			14'd6211: ff_rdata <= 8'hF5;
			14'd6212: ff_rdata <= 8'h01;
			14'd6213: ff_rdata <= 8'h25;
			14'd6214: ff_rdata <= 8'h00;
			14'd6215: ff_rdata <= 8'hED;
			14'd6216: ff_rdata <= 8'hB0;
			14'd6217: ff_rdata <= 8'hE1;
			14'd6218: ff_rdata <= 8'hCD;
			14'd6219: ff_rdata <= 8'hB5;
			14'd6220: ff_rdata <= 8'h67;
			14'd6221: ff_rdata <= 8'hE3;
			14'd6222: ff_rdata <= 8'hE5;
			14'd6223: ff_rdata <= 8'hCD;
			14'd6224: ff_rdata <= 8'hD3;
			14'd6225: ff_rdata <= 8'h67;
			14'd6226: ff_rdata <= 8'hCD;
			14'd6227: ff_rdata <= 8'h34;
			14'd6228: ff_rdata <= 8'h68;
			14'd6229: ff_rdata <= 8'h7B;
			14'd6230: ff_rdata <= 8'hB7;
			14'd6231: ff_rdata <= 8'h20;
			14'd6232: ff_rdata <= 8'h05;
			14'd6233: ff_rdata <= 8'h11;
			14'd6234: ff_rdata <= 8'h01;
			14'd6235: ff_rdata <= 8'hA0;
			14'd6236: ff_rdata <= 8'h0E;
			14'd6237: ff_rdata <= 8'h57;
			14'd6238: ff_rdata <= 8'hF1;
			14'd6239: ff_rdata <= 8'hF5;
			14'd6240: ff_rdata <= 8'hCD;
			14'd6241: ff_rdata <= 8'h02;
			14'd6242: ff_rdata <= 8'h5F;
			14'd6243: ff_rdata <= 8'hAF;
			14'd6244: ff_rdata <= 8'hDD;
			14'd6245: ff_rdata <= 8'h77;
			14'd6246: ff_rdata <= 8'h00;
			14'd6247: ff_rdata <= 8'hF1;
			14'd6248: ff_rdata <= 8'hF5;
			14'd6249: ff_rdata <= 8'hCD;
			14'd6250: ff_rdata <= 8'hE0;
			14'd6251: ff_rdata <= 8'h67;
			14'd6252: ff_rdata <= 8'h73;
			14'd6253: ff_rdata <= 8'h23;
			14'd6254: ff_rdata <= 8'h72;
			14'd6255: ff_rdata <= 8'h23;
			14'd6256: ff_rdata <= 8'h71;
			14'd6257: ff_rdata <= 8'h23;
			14'd6258: ff_rdata <= 8'h54;
			14'd6259: ff_rdata <= 8'h5D;
			14'd6260: ff_rdata <= 8'h01;
			14'd6261: ff_rdata <= 8'h1C;
			14'd6262: ff_rdata <= 8'h00;
			14'd6263: ff_rdata <= 8'h09;
			14'd6264: ff_rdata <= 8'hEB;
			14'd6265: ff_rdata <= 8'h73;
			14'd6266: ff_rdata <= 8'h23;
			14'd6267: ff_rdata <= 8'h72;
			14'd6268: ff_rdata <= 8'hC1;
			14'd6269: ff_rdata <= 8'hE1;
			14'd6270: ff_rdata <= 8'h04;
			14'd6271: ff_rdata <= 8'h3A;
			14'd6272: ff_rdata <= 8'h91;
			14'd6273: ff_rdata <= 8'hF9;
			14'd6274: ff_rdata <= 8'h3D;
			14'd6275: ff_rdata <= 8'hB8;
			14'd6276: ff_rdata <= 8'h38;
			14'd6277: ff_rdata <= 8'h22;
			14'd6278: ff_rdata <= 8'h2B;
			14'd6279: ff_rdata <= 8'hCD;
			14'd6280: ff_rdata <= 8'hAF;
			14'd6281: ff_rdata <= 8'h67;
			14'd6282: ff_rdata <= 8'h28;
			14'd6283: ff_rdata <= 8'h06;
			14'd6284: ff_rdata <= 8'hC5;
			14'd6285: ff_rdata <= 8'hCD;
			14'd6286: ff_rdata <= 8'hDF;
			14'd6287: ff_rdata <= 8'h55;
			14'd6288: ff_rdata <= 8'h18;
			14'd6289: ff_rdata <= 8'hAB;
			14'd6290: ff_rdata <= 8'h78;
			14'd6291: ff_rdata <= 8'h32;
			14'd6292: ff_rdata <= 8'h38;
			14'd6293: ff_rdata <= 8'hFB;
			14'd6294: ff_rdata <= 8'hC5;
			14'd6295: ff_rdata <= 8'hE5;
			14'd6296: ff_rdata <= 8'hCD;
			14'd6297: ff_rdata <= 8'hAF;
			14'd6298: ff_rdata <= 8'h59;
			14'd6299: ff_rdata <= 8'hE1;
			14'd6300: ff_rdata <= 8'hC1;
			14'd6301: ff_rdata <= 8'hCD;
			14'd6302: ff_rdata <= 8'h95;
			14'd6303: ff_rdata <= 8'h59;
			14'd6304: ff_rdata <= 8'h04;
			14'd6305: ff_rdata <= 8'h3A;
			14'd6306: ff_rdata <= 8'h91;
			14'd6307: ff_rdata <= 8'hF9;
			14'd6308: ff_rdata <= 8'h3D;
			14'd6309: ff_rdata <= 8'hB8;
			14'd6310: ff_rdata <= 8'h30;
			14'd6311: ff_rdata <= 8'hEA;
			14'd6312: ff_rdata <= 8'h2B;
			14'd6313: ff_rdata <= 8'hCD;
			14'd6314: ff_rdata <= 8'hAF;
			14'd6315: ff_rdata <= 8'h67;
			14'd6316: ff_rdata <= 8'hC2;
			14'd6317: ff_rdata <= 8'h6D;
			14'd6318: ff_rdata <= 8'h67;
			14'd6319: ff_rdata <= 8'hE5;
			14'd6320: ff_rdata <= 8'hAF;
			14'd6321: ff_rdata <= 8'hF5;
			14'd6322: ff_rdata <= 8'h32;
			14'd6323: ff_rdata <= 8'h38;
			14'd6324: ff_rdata <= 8'hFB;
			14'd6325: ff_rdata <= 8'h4F;
			14'd6326: ff_rdata <= 8'h3A;
			14'd6327: ff_rdata <= 8'h91;
			14'd6328: ff_rdata <= 8'hF9;
			14'd6329: ff_rdata <= 8'h91;
			14'd6330: ff_rdata <= 8'hD6;
			14'd6331: ff_rdata <= 8'h04;
			14'd6332: ff_rdata <= 8'h21;
			14'd6333: ff_rdata <= 8'hE2;
			14'd6334: ff_rdata <= 8'h59;
			14'd6335: ff_rdata <= 8'h38;
			14'd6336: ff_rdata <= 8'h0F;
			14'd6337: ff_rdata <= 8'h21;
			14'd6338: ff_rdata <= 8'h70;
			14'd6339: ff_rdata <= 8'h5C;
			14'd6340: ff_rdata <= 8'h20;
			14'd6341: ff_rdata <= 8'h0A;
			14'd6342: ff_rdata <= 8'h3A;
			14'd6343: ff_rdata <= 8'h8E;
			14'd6344: ff_rdata <= 8'hF9;
			14'd6345: ff_rdata <= 8'hE6;
			14'd6346: ff_rdata <= 8'h01;
			14'd6347: ff_rdata <= 8'h28;
			14'd6348: ff_rdata <= 8'h03;
			14'd6349: ff_rdata <= 8'h21;
			14'd6350: ff_rdata <= 8'hA2;
			14'd6351: ff_rdata <= 8'h5F;
			14'd6352: ff_rdata <= 8'h22;
			14'd6353: ff_rdata <= 8'h56;
			14'd6354: ff_rdata <= 8'hF9;
			14'd6355: ff_rdata <= 8'h79;
			14'd6356: ff_rdata <= 8'h47;
			14'd6357: ff_rdata <= 8'hCD;
			14'd6358: ff_rdata <= 8'hD5;
			14'd6359: ff_rdata <= 8'h59;
			14'd6360: ff_rdata <= 8'hDA;
			14'd6361: ff_rdata <= 8'h57;
			14'd6362: ff_rdata <= 8'h59;
			14'd6363: ff_rdata <= 8'h78;
			14'd6364: ff_rdata <= 8'hCD;
			14'd6365: ff_rdata <= 8'hE0;
			14'd6366: ff_rdata <= 8'h67;
			14'd6367: ff_rdata <= 8'h7E;
			14'd6368: ff_rdata <= 8'hB7;
			14'd6369: ff_rdata <= 8'hCA;
			14'd6370: ff_rdata <= 8'h57;
			14'd6371: ff_rdata <= 8'h59;
			14'd6372: ff_rdata <= 8'h32;
			14'd6373: ff_rdata <= 8'h3B;
			14'd6374: ff_rdata <= 8'hFB;
			14'd6375: ff_rdata <= 8'h23;
			14'd6376: ff_rdata <= 8'h5E;
			14'd6377: ff_rdata <= 8'h23;
			14'd6378: ff_rdata <= 8'h56;
			14'd6379: ff_rdata <= 8'h23;
			14'd6380: ff_rdata <= 8'hED;
			14'd6381: ff_rdata <= 8'h53;
			14'd6382: ff_rdata <= 8'h3C;
			14'd6383: ff_rdata <= 8'hFB;
			14'd6384: ff_rdata <= 8'h5E;
			14'd6385: ff_rdata <= 8'h23;
			14'd6386: ff_rdata <= 8'h56;
			14'd6387: ff_rdata <= 8'h23;
			14'd6388: ff_rdata <= 8'hE5;
			14'd6389: ff_rdata <= 8'h2E;
			14'd6390: ff_rdata <= 8'h24;
			14'd6391: ff_rdata <= 8'hCD;
			14'd6392: ff_rdata <= 8'hE4;
			14'd6393: ff_rdata <= 8'h67;
			14'd6394: ff_rdata <= 8'hE5;
			14'd6395: ff_rdata <= 8'h2A;
			14'd6396: ff_rdata <= 8'h36;
			14'd6397: ff_rdata <= 8'hFB;
			14'd6398: ff_rdata <= 8'h2B;
			14'd6399: ff_rdata <= 8'hC1;
			14'd6400: ff_rdata <= 8'hF3;
			14'd6401: ff_rdata <= 8'hCD;
			14'd6402: ff_rdata <= 8'h27;
			14'd6403: ff_rdata <= 8'h68;
			14'd6404: ff_rdata <= 8'hD1;
			14'd6405: ff_rdata <= 8'h60;
			14'd6406: ff_rdata <= 8'h69;
			14'd6407: ff_rdata <= 8'hF9;
			14'd6408: ff_rdata <= 8'hFB;
			14'd6409: ff_rdata <= 8'hCD;
			14'd6410: ff_rdata <= 8'hAF;
			14'd6411: ff_rdata <= 8'h59;
			14'd6412: ff_rdata <= 8'hC3;
			14'd6413: ff_rdata <= 8'hC6;
			14'd6414: ff_rdata <= 8'h65;
			14'd6415: ff_rdata <= 8'h3A;
			14'd6416: ff_rdata <= 8'h3B;
			14'd6417: ff_rdata <= 8'hFB;
			14'd6418: ff_rdata <= 8'hB7;
			14'd6419: ff_rdata <= 8'h20;
			14'd6420: ff_rdata <= 8'h03;
			14'd6421: ff_rdata <= 8'hCD;
			14'd6422: ff_rdata <= 8'h95;
			14'd6423: ff_rdata <= 8'h59;
			14'd6424: ff_rdata <= 8'h3A;
			14'd6425: ff_rdata <= 8'h38;
			14'd6426: ff_rdata <= 8'hFB;
			14'd6427: ff_rdata <= 8'hCD;
			14'd6428: ff_rdata <= 8'hE0;
			14'd6429: ff_rdata <= 8'h67;
			14'd6430: ff_rdata <= 8'h3A;
			14'd6431: ff_rdata <= 8'h3B;
			14'd6432: ff_rdata <= 8'hFB;
			14'd6433: ff_rdata <= 8'h77;
			14'd6434: ff_rdata <= 8'h23;
			14'd6435: ff_rdata <= 8'hED;
			14'd6436: ff_rdata <= 8'h5B;
			14'd6437: ff_rdata <= 8'h3C;
			14'd6438: ff_rdata <= 8'hFB;
			14'd6439: ff_rdata <= 8'h73;
			14'd6440: ff_rdata <= 8'h23;
			14'd6441: ff_rdata <= 8'h72;
			14'd6442: ff_rdata <= 8'h21;
			14'd6443: ff_rdata <= 8'h00;
			14'd6444: ff_rdata <= 8'h00;
			14'd6445: ff_rdata <= 8'h39;
			14'd6446: ff_rdata <= 8'hEB;
			14'd6447: ff_rdata <= 8'h2A;
			14'd6448: ff_rdata <= 8'h36;
			14'd6449: ff_rdata <= 8'hFB;
			14'd6450: ff_rdata <= 8'hF3;
			14'd6451: ff_rdata <= 8'hF9;
			14'd6452: ff_rdata <= 8'hC1;
			14'd6453: ff_rdata <= 8'hC1;
			14'd6454: ff_rdata <= 8'hC1;
			14'd6455: ff_rdata <= 8'hE5;
			14'd6456: ff_rdata <= 8'hB7;
			14'd6457: ff_rdata <= 8'hED;
			14'd6458: ff_rdata <= 8'h52;
			14'd6459: ff_rdata <= 8'h28;
			14'd6460: ff_rdata <= 8'h18;
			14'd6461: ff_rdata <= 8'h3E;
			14'd6462: ff_rdata <= 8'hF0;
			14'd6463: ff_rdata <= 8'hA5;
			14'd6464: ff_rdata <= 8'hB4;
			14'd6465: ff_rdata <= 8'hC2;
			14'd6466: ff_rdata <= 8'h70;
			14'd6467: ff_rdata <= 8'h67;
			14'd6468: ff_rdata <= 8'h2E;
			14'd6469: ff_rdata <= 8'h24;
			14'd6470: ff_rdata <= 8'hCD;
			14'd6471: ff_rdata <= 8'hE4;
			14'd6472: ff_rdata <= 8'h67;
			14'd6473: ff_rdata <= 8'hC1;
			14'd6474: ff_rdata <= 8'h0B;
			14'd6475: ff_rdata <= 8'hCD;
			14'd6476: ff_rdata <= 8'h27;
			14'd6477: ff_rdata <= 8'h68;
			14'd6478: ff_rdata <= 8'hE1;
			14'd6479: ff_rdata <= 8'h2B;
			14'd6480: ff_rdata <= 8'h70;
			14'd6481: ff_rdata <= 8'h2B;
			14'd6482: ff_rdata <= 8'h71;
			14'd6483: ff_rdata <= 8'h18;
			14'd6484: ff_rdata <= 8'h02;
			14'd6485: ff_rdata <= 8'hC1;
			14'd6486: ff_rdata <= 8'hC1;
			14'd6487: ff_rdata <= 8'hFB;
			14'd6488: ff_rdata <= 8'hF1;
			14'd6489: ff_rdata <= 8'h3C;
			14'd6490: ff_rdata <= 8'h21;
			14'd6491: ff_rdata <= 8'h91;
			14'd6492: ff_rdata <= 8'hF9;
			14'd6493: ff_rdata <= 8'hBE;
			14'd6494: ff_rdata <= 8'hDA;
			14'd6495: ff_rdata <= 8'hB1;
			14'd6496: ff_rdata <= 8'h58;
			14'd6497: ff_rdata <= 8'hF3;
			14'd6498: ff_rdata <= 8'hCD;
			14'd6499: ff_rdata <= 8'hB1;
			14'd6500: ff_rdata <= 8'h63;
			14'd6501: ff_rdata <= 8'h28;
			14'd6502: ff_rdata <= 8'h28;
			14'd6503: ff_rdata <= 8'h3A;
			14'd6504: ff_rdata <= 8'h35;
			14'd6505: ff_rdata <= 8'hFB;
			14'd6506: ff_rdata <= 8'h07;
			14'd6507: ff_rdata <= 8'h38;
			14'd6508: ff_rdata <= 8'h0B;
			14'd6509: ff_rdata <= 8'h21;
			14'd6510: ff_rdata <= 8'h97;
			14'd6511: ff_rdata <= 8'hF9;
			14'd6512: ff_rdata <= 8'h34;
			14'd6513: ff_rdata <= 8'h7E;
			14'd6514: ff_rdata <= 8'h32;
			14'd6515: ff_rdata <= 8'h40;
			14'd6516: ff_rdata <= 8'hFB;
			14'd6517: ff_rdata <= 8'hCD;
			14'd6518: ff_rdata <= 8'h3D;
			14'd6519: ff_rdata <= 8'h68;
			14'd6520: ff_rdata <= 8'hFB;
			14'd6521: ff_rdata <= 8'h21;
			14'd6522: ff_rdata <= 8'h35;
			14'd6523: ff_rdata <= 8'hFB;
			14'd6524: ff_rdata <= 8'hCB;
			14'd6525: ff_rdata <= 8'hFE;
			14'd6526: ff_rdata <= 8'h7E;
			14'd6527: ff_rdata <= 8'h21;
			14'd6528: ff_rdata <= 8'h93;
			14'd6529: ff_rdata <= 8'hF9;
			14'd6530: ff_rdata <= 8'hBE;
			14'd6531: ff_rdata <= 8'hC2;
			14'd6532: ff_rdata <= 8'hB0;
			14'd6533: ff_rdata <= 8'h58;
			14'd6534: ff_rdata <= 8'h3A;
			14'd6535: ff_rdata <= 8'h98;
			14'd6536: ff_rdata <= 8'hF9;
			14'd6537: ff_rdata <= 8'hB7;
			14'd6538: ff_rdata <= 8'hC4;
			14'd6539: ff_rdata <= 8'h9D;
			14'd6540: ff_rdata <= 8'h63;
			14'd6541: ff_rdata <= 8'h30;
			14'd6542: ff_rdata <= 8'h04;
			14'd6543: ff_rdata <= 8'hCD;
			14'd6544: ff_rdata <= 8'h8D;
			14'd6545: ff_rdata <= 8'h65;
			14'd6546: ff_rdata <= 8'hFB;
			14'd6547: ff_rdata <= 8'hE1;
			14'd6548: ff_rdata <= 8'hC9;
			14'd6549: ff_rdata <= 8'h3A;
			14'd6550: ff_rdata <= 8'h35;
			14'd6551: ff_rdata <= 8'hFB;
			14'd6552: ff_rdata <= 8'h3C;
			14'd6553: ff_rdata <= 8'h32;
			14'd6554: ff_rdata <= 8'h35;
			14'd6555: ff_rdata <= 8'hFB;
			14'd6556: ff_rdata <= 8'h1E;
			14'd6557: ff_rdata <= 8'hFF;
			14'd6558: ff_rdata <= 8'hE5;
			14'd6559: ff_rdata <= 8'hC5;
			14'd6560: ff_rdata <= 8'hD5;
			14'd6561: ff_rdata <= 8'h3A;
			14'd6562: ff_rdata <= 8'h38;
			14'd6563: ff_rdata <= 8'hFB;
			14'd6564: ff_rdata <= 8'hF3;
			14'd6565: ff_rdata <= 8'hCD;
			14'd6566: ff_rdata <= 8'hF9;
			14'd6567: ff_rdata <= 8'h66;
			14'd6568: ff_rdata <= 8'hFB;
			14'd6569: ff_rdata <= 8'hD1;
			14'd6570: ff_rdata <= 8'h28;
			14'd6571: ff_rdata <= 8'hF4;
			14'd6572: ff_rdata <= 8'hC1;
			14'd6573: ff_rdata <= 8'hE1;
			14'd6574: ff_rdata <= 8'hC9;
			14'd6575: ff_rdata <= 8'h21;
			14'd6576: ff_rdata <= 8'h38;
			14'd6577: ff_rdata <= 8'hFB;
			14'd6578: ff_rdata <= 8'h3A;
			14'd6579: ff_rdata <= 8'h92;
			14'd6580: ff_rdata <= 8'hF9;
			14'd6581: ff_rdata <= 8'h3D;
			14'd6582: ff_rdata <= 8'hBE;
			14'd6583: ff_rdata <= 8'hC0;
			14'd6584: ff_rdata <= 8'h3A;
			14'd6585: ff_rdata <= 8'h7F;
			14'd6586: ff_rdata <= 8'hF9;
			14'd6587: ff_rdata <= 8'h21;
			14'd6588: ff_rdata <= 8'h80;
			14'd6589: ff_rdata <= 8'hF9;
			14'd6590: ff_rdata <= 8'hBE;
			14'd6591: ff_rdata <= 8'hC8;
			14'd6592: ff_rdata <= 8'h77;
			14'd6593: ff_rdata <= 8'h3E;
			14'd6594: ff_rdata <= 8'h88;
			14'd6595: ff_rdata <= 8'hB6;
			14'd6596: ff_rdata <= 8'h5F;
			14'd6597: ff_rdata <= 8'hE5;
			14'd6598: ff_rdata <= 8'hC5;
			14'd6599: ff_rdata <= 8'hD5;
			14'd6600: ff_rdata <= 8'h3A;
			14'd6601: ff_rdata <= 8'h38;
			14'd6602: ff_rdata <= 8'hFB;
			14'd6603: ff_rdata <= 8'hF3;
			14'd6604: ff_rdata <= 8'hCD;
			14'd6605: ff_rdata <= 8'hF9;
			14'd6606: ff_rdata <= 8'h66;
			14'd6607: ff_rdata <= 8'hD1;
			14'd6608: ff_rdata <= 8'h20;
			14'd6609: ff_rdata <= 8'hDA;
			14'd6610: ff_rdata <= 8'hFB;
			14'd6611: ff_rdata <= 8'h18;
			14'd6612: ff_rdata <= 8'hF2;
			14'd6613: ff_rdata <= 8'h3A;
			14'd6614: ff_rdata <= 8'h38;
			14'd6615: ff_rdata <= 8'hFB;
			14'd6616: ff_rdata <= 8'hC5;
			14'd6617: ff_rdata <= 8'hF3;
			14'd6618: ff_rdata <= 8'hCD;
			14'd6619: ff_rdata <= 8'h41;
			14'd6620: ff_rdata <= 8'h67;
			14'd6621: ff_rdata <= 8'hFB;
			14'd6622: ff_rdata <= 8'hC1;
			14'd6623: ff_rdata <= 8'hFE;
			14'd6624: ff_rdata <= 8'h08;
			14'd6625: ff_rdata <= 8'hC9;
			14'd6626: ff_rdata <= 8'h41;
			14'd6627: ff_rdata <= 8'h1D;
			14'd6628: ff_rdata <= 8'h5B;
			14'd6629: ff_rdata <= 8'hCD;
			14'd6630: ff_rdata <= 8'h54;
			14'd6631: ff_rdata <= 8'h5A;
			14'd6632: ff_rdata <= 8'hD6;
			14'd6633: ff_rdata <= 8'h3D;
			14'd6634: ff_rdata <= 8'h5A;
			14'd6635: ff_rdata <= 8'hD3;
			14'd6636: ff_rdata <= 8'h76;
			14'd6637: ff_rdata <= 8'h5A;
			14'd6638: ff_rdata <= 8'hCE;
			14'd6639: ff_rdata <= 8'hDA;
			14'd6640: ff_rdata <= 8'h5A;
			14'd6641: ff_rdata <= 8'hCF;
			14'd6642: ff_rdata <= 8'hA6;
			14'd6643: ff_rdata <= 8'h5A;
			14'd6644: ff_rdata <= 8'hD2;
			14'd6645: ff_rdata <= 8'hB5;
			14'd6646: ff_rdata <= 8'h5A;
			14'd6647: ff_rdata <= 8'hD4;
			14'd6648: ff_rdata <= 8'h99;
			14'd6649: ff_rdata <= 8'h5A;
			14'd6650: ff_rdata <= 8'hCC;
			14'd6651: ff_rdata <= 8'h80;
			14'd6652: ff_rdata <= 8'h5A;
			14'd6653: ff_rdata <= 8'h58;
			14'd6654: ff_rdata <= 8'hDB;
			14'd6655: ff_rdata <= 8'h66;
			14'd6656: ff_rdata <= 8'h3E;
			14'd6657: ff_rdata <= 8'hAB;
			14'd6658: ff_rdata <= 8'h5D;
			14'd6659: ff_rdata <= 8'h3C;
			14'd6660: ff_rdata <= 8'hB8;
			14'd6661: ff_rdata <= 8'h5D;
			14'd6662: ff_rdata <= 8'hD9;
			14'd6663: ff_rdata <= 8'h04;
			14'd6664: ff_rdata <= 8'h5C;
			14'd6665: ff_rdata <= 8'hD1;
			14'd6666: ff_rdata <= 8'h1A;
			14'd6667: ff_rdata <= 8'h5C;
			14'd6668: ff_rdata <= 8'h40;
			14'd6669: ff_rdata <= 8'h29;
			14'd6670: ff_rdata <= 8'h5C;
			14'd6671: ff_rdata <= 8'h26;
			14'd6672: ff_rdata <= 8'h03;
			14'd6673: ff_rdata <= 8'h5C;
			14'd6674: ff_rdata <= 8'hDA;
			14'd6675: ff_rdata <= 8'h25;
			14'd6676: ff_rdata <= 8'h5C;
			14'd6677: ff_rdata <= 8'h00;
			14'd6678: ff_rdata <= 8'h10;
			14'd6679: ff_rdata <= 8'h12;
			14'd6680: ff_rdata <= 8'h14;
			14'd6681: ff_rdata <= 8'h16;
			14'd6682: ff_rdata <= 8'h00;
			14'd6683: ff_rdata <= 8'h00;
			14'd6684: ff_rdata <= 8'h02;
			14'd6685: ff_rdata <= 8'h04;
			14'd6686: ff_rdata <= 8'h06;
			14'd6687: ff_rdata <= 8'h08;
			14'd6688: ff_rdata <= 8'h0A;
			14'd6689: ff_rdata <= 8'h0A;
			14'd6690: ff_rdata <= 8'h0C;
			14'd6691: ff_rdata <= 8'h0E;
			14'd6692: ff_rdata <= 8'h10;
			14'd6693: ff_rdata <= 8'h5D;
			14'd6694: ff_rdata <= 8'h0D;
			14'd6695: ff_rdata <= 8'h9C;
			14'd6696: ff_rdata <= 8'h0C;
			14'd6697: ff_rdata <= 8'hE7;
			14'd6698: ff_rdata <= 8'h0B;
			14'd6699: ff_rdata <= 8'h3C;
			14'd6700: ff_rdata <= 8'h0B;
			14'd6701: ff_rdata <= 8'h9B;
			14'd6702: ff_rdata <= 8'h0A;
			14'd6703: ff_rdata <= 8'h02;
			14'd6704: ff_rdata <= 8'h0A;
			14'd6705: ff_rdata <= 8'h73;
			14'd6706: ff_rdata <= 8'h09;
			14'd6707: ff_rdata <= 8'hEB;
			14'd6708: ff_rdata <= 8'h08;
			14'd6709: ff_rdata <= 8'h6B;
			14'd6710: ff_rdata <= 8'h08;
			14'd6711: ff_rdata <= 8'hF2;
			14'd6712: ff_rdata <= 8'h07;
			14'd6713: ff_rdata <= 8'h80;
			14'd6714: ff_rdata <= 8'h07;
			14'd6715: ff_rdata <= 8'h14;
			14'd6716: ff_rdata <= 8'h07;
			14'd6717: ff_rdata <= 8'h38;
			14'd6718: ff_rdata <= 8'h02;
			14'd6719: ff_rdata <= 8'h1E;
			14'd6720: ff_rdata <= 8'h08;
			14'd6721: ff_rdata <= 8'h3E;
			14'd6722: ff_rdata <= 8'h0F;
			14'd6723: ff_rdata <= 8'hBB;
			14'd6724: ff_rdata <= 8'h38;
			14'd6725: ff_rdata <= 8'h50;
			14'd6726: ff_rdata <= 8'hCD;
			14'd6727: ff_rdata <= 8'h41;
			14'd6728: ff_rdata <= 8'h5C;
			14'd6729: ff_rdata <= 8'h2E;
			14'd6730: ff_rdata <= 8'h12;
			14'd6731: ff_rdata <= 8'hCD;
			14'd6732: ff_rdata <= 8'hE4;
			14'd6733: ff_rdata <= 8'h67;
			14'd6734: ff_rdata <= 8'h3E;
			14'd6735: ff_rdata <= 8'h40;
			14'd6736: ff_rdata <= 8'hA6;
			14'd6737: ff_rdata <= 8'hB3;
			14'd6738: ff_rdata <= 8'h77;
			14'd6739: ff_rdata <= 8'hC9;
			14'd6740: ff_rdata <= 8'h7B;
			14'd6741: ff_rdata <= 8'h38;
			14'd6742: ff_rdata <= 8'h03;
			14'd6743: ff_rdata <= 8'h2F;
			14'd6744: ff_rdata <= 8'h3C;
			14'd6745: ff_rdata <= 8'h5F;
			14'd6746: ff_rdata <= 8'hB2;
			14'd6747: ff_rdata <= 8'h28;
			14'd6748: ff_rdata <= 8'h39;
			14'd6749: ff_rdata <= 8'h2E;
			14'd6750: ff_rdata <= 8'h13;
			14'd6751: ff_rdata <= 8'hCD;
			14'd6752: ff_rdata <= 8'hE4;
			14'd6753: ff_rdata <= 8'h67;
			14'd6754: ff_rdata <= 8'hE5;
			14'd6755: ff_rdata <= 8'h7E;
			14'd6756: ff_rdata <= 8'h23;
			14'd6757: ff_rdata <= 8'h66;
			14'd6758: ff_rdata <= 8'h6F;
			14'd6759: ff_rdata <= 8'hCD;
			14'd6760: ff_rdata <= 8'hD4;
			14'd6761: ff_rdata <= 8'h68;
			14'd6762: ff_rdata <= 8'hE1;
			14'd6763: ff_rdata <= 8'hC8;
			14'd6764: ff_rdata <= 8'h73;
			14'd6765: ff_rdata <= 8'h23;
			14'd6766: ff_rdata <= 8'h72;
			14'd6767: ff_rdata <= 8'h2B;
			14'd6768: ff_rdata <= 8'h2B;
			14'd6769: ff_rdata <= 8'h3E;
			14'd6770: ff_rdata <= 8'h40;
			14'd6771: ff_rdata <= 8'hB6;
			14'd6772: ff_rdata <= 8'h77;
			14'd6773: ff_rdata <= 8'hC9;
			14'd6774: ff_rdata <= 8'h7B;
			14'd6775: ff_rdata <= 8'hFE;
			14'd6776: ff_rdata <= 8'h10;
			14'd6777: ff_rdata <= 8'h30;
			14'd6778: ff_rdata <= 8'h1B;
			14'd6779: ff_rdata <= 8'hF6;
			14'd6780: ff_rdata <= 8'h10;
			14'd6781: ff_rdata <= 8'h5F;
			14'd6782: ff_rdata <= 8'h18;
			14'd6783: ff_rdata <= 8'hC6;
			14'd6784: ff_rdata <= 8'h38;
			14'd6785: ff_rdata <= 8'h02;
			14'd6786: ff_rdata <= 8'h1E;
			14'd6787: ff_rdata <= 8'h04;
			14'd6788: ff_rdata <= 8'h7B;
			14'd6789: ff_rdata <= 8'hFE;
			14'd6790: ff_rdata <= 8'h41;
			14'd6791: ff_rdata <= 8'h30;
			14'd6792: ff_rdata <= 8'h0D;
			14'd6793: ff_rdata <= 8'h2E;
			14'd6794: ff_rdata <= 8'h10;
			14'd6795: ff_rdata <= 8'hCD;
			14'd6796: ff_rdata <= 8'hE4;
			14'd6797: ff_rdata <= 8'h67;
			14'd6798: ff_rdata <= 8'hCD;
			14'd6799: ff_rdata <= 8'h41;
			14'd6800: ff_rdata <= 8'h5C;
			14'd6801: ff_rdata <= 8'hB3;
			14'd6802: ff_rdata <= 8'h28;
			14'd6803: ff_rdata <= 8'h02;
			14'd6804: ff_rdata <= 8'h77;
			14'd6805: ff_rdata <= 8'hC9;
			14'd6806: ff_rdata <= 8'hC3;
			14'd6807: ff_rdata <= 8'h70;
			14'd6808: ff_rdata <= 8'h67;
			14'd6809: ff_rdata <= 8'h38;
			14'd6810: ff_rdata <= 8'h02;
			14'd6811: ff_rdata <= 8'h1E;
			14'd6812: ff_rdata <= 8'h78;
			14'd6813: ff_rdata <= 8'h7B;
			14'd6814: ff_rdata <= 8'hFE;
			14'd6815: ff_rdata <= 8'h20;
			14'd6816: ff_rdata <= 8'h38;
			14'd6817: ff_rdata <= 8'hF4;
			14'd6818: ff_rdata <= 8'h2E;
			14'd6819: ff_rdata <= 8'h11;
			14'd6820: ff_rdata <= 8'h18;
			14'd6821: ff_rdata <= 8'hE5;
			14'd6822: ff_rdata <= 8'h38;
			14'd6823: ff_rdata <= 8'h02;
			14'd6824: ff_rdata <= 8'h1E;
			14'd6825: ff_rdata <= 8'h04;
			14'd6826: ff_rdata <= 8'h7B;
			14'd6827: ff_rdata <= 8'hFE;
			14'd6828: ff_rdata <= 8'h09;
			14'd6829: ff_rdata <= 8'h30;
			14'd6830: ff_rdata <= 8'hE7;
			14'd6831: ff_rdata <= 8'h2E;
			14'd6832: ff_rdata <= 8'h0F;
			14'd6833: ff_rdata <= 8'h18;
			14'd6834: ff_rdata <= 8'hD8;
			14'd6835: ff_rdata <= 8'hAF;
			14'd6836: ff_rdata <= 8'h57;
			14'd6837: ff_rdata <= 8'h38;
			14'd6838: ff_rdata <= 8'h02;
			14'd6839: ff_rdata <= 8'h1E;
			14'd6840: ff_rdata <= 8'h04;
			14'd6841: ff_rdata <= 8'hAF;
			14'd6842: ff_rdata <= 8'hB2;
			14'd6843: ff_rdata <= 8'h20;
			14'd6844: ff_rdata <= 8'hD9;
			14'd6845: ff_rdata <= 8'hB3;
			14'd6846: ff_rdata <= 8'h28;
			14'd6847: ff_rdata <= 8'hD6;
			14'd6848: ff_rdata <= 8'hFE;
			14'd6849: ff_rdata <= 8'h41;
			14'd6850: ff_rdata <= 8'h30;
			14'd6851: ff_rdata <= 8'hD2;
			14'd6852: ff_rdata <= 8'h21;
			14'd6853: ff_rdata <= 8'h00;
			14'd6854: ff_rdata <= 8'h00;
			14'd6855: ff_rdata <= 8'hE5;
			14'd6856: ff_rdata <= 8'h2E;
			14'd6857: ff_rdata <= 8'h10;
			14'd6858: ff_rdata <= 8'hCD;
			14'd6859: ff_rdata <= 8'hE4;
			14'd6860: ff_rdata <= 8'h67;
			14'd6861: ff_rdata <= 8'hE5;
			14'd6862: ff_rdata <= 8'h23;
			14'd6863: ff_rdata <= 8'h23;
			14'd6864: ff_rdata <= 8'h7E;
			14'd6865: ff_rdata <= 8'h32;
			14'd6866: ff_rdata <= 8'h39;
			14'd6867: ff_rdata <= 8'hFB;
			14'd6868: ff_rdata <= 8'h36;
			14'd6869: ff_rdata <= 8'h80;
			14'd6870: ff_rdata <= 8'h2B;
			14'd6871: ff_rdata <= 8'h2B;
			14'd6872: ff_rdata <= 8'h18;
			14'd6873: ff_rdata <= 8'h7E;
			14'd6874: ff_rdata <= 8'h30;
			14'd6875: ff_rdata <= 8'hBA;
			14'd6876: ff_rdata <= 8'hCD;
			14'd6877: ff_rdata <= 8'h41;
			14'd6878: ff_rdata <= 8'h5C;
			14'd6879: ff_rdata <= 8'hB3;
			14'd6880: ff_rdata <= 8'h28;
			14'd6881: ff_rdata <= 8'hE2;
			14'd6882: ff_rdata <= 8'hFE;
			14'd6883: ff_rdata <= 8'h61;
			14'd6884: ff_rdata <= 8'h30;
			14'd6885: ff_rdata <= 8'hB0;
			14'd6886: ff_rdata <= 8'h7B;
			14'd6887: ff_rdata <= 8'h06;
			14'd6888: ff_rdata <= 8'h00;
			14'd6889: ff_rdata <= 8'h58;
			14'd6890: ff_rdata <= 8'hD6;
			14'd6891: ff_rdata <= 8'h0C;
			14'd6892: ff_rdata <= 8'h1C;
			14'd6893: ff_rdata <= 8'h30;
			14'd6894: ff_rdata <= 8'hFB;
			14'd6895: ff_rdata <= 8'hC6;
			14'd6896: ff_rdata <= 8'h0C;
			14'd6897: ff_rdata <= 8'h87;
			14'd6898: ff_rdata <= 8'h4F;
			14'd6899: ff_rdata <= 8'hC3;
			14'd6900: ff_rdata <= 8'h2D;
			14'd6901: ff_rdata <= 8'h5B;
			14'd6902: ff_rdata <= 8'h41;
			14'd6903: ff_rdata <= 8'h79;
			14'd6904: ff_rdata <= 8'hD6;
			14'd6905: ff_rdata <= 8'h40;
			14'd6906: ff_rdata <= 8'h87;
			14'd6907: ff_rdata <= 8'h4F;
			14'd6908: ff_rdata <= 8'hCD;
			14'd6909: ff_rdata <= 8'h1A;
			14'd6910: ff_rdata <= 8'h66;
			14'd6911: ff_rdata <= 8'h28;
			14'd6912: ff_rdata <= 8'h1A;
			14'd6913: ff_rdata <= 8'hFE;
			14'd6914: ff_rdata <= 8'h23;
			14'd6915: ff_rdata <= 8'hC8;
			14'd6916: ff_rdata <= 8'hFE;
			14'd6917: ff_rdata <= 8'h2B;
			14'd6918: ff_rdata <= 8'hC8;
			14'd6919: ff_rdata <= 8'hFE;
			14'd6920: ff_rdata <= 8'h2D;
			14'd6921: ff_rdata <= 8'h28;
			14'd6922: ff_rdata <= 8'h05;
			14'd6923: ff_rdata <= 8'hCD;
			14'd6924: ff_rdata <= 8'h40;
			14'd6925: ff_rdata <= 8'h66;
			14'd6926: ff_rdata <= 8'h18;
			14'd6927: ff_rdata <= 8'h0B;
			14'd6928: ff_rdata <= 8'h0D;
			14'd6929: ff_rdata <= 8'h78;
			14'd6930: ff_rdata <= 8'hFE;
			14'd6931: ff_rdata <= 8'h43;
			14'd6932: ff_rdata <= 8'h28;
			14'd6933: ff_rdata <= 8'h04;
			14'd6934: ff_rdata <= 8'hFE;
			14'd6935: ff_rdata <= 8'h46;
			14'd6936: ff_rdata <= 8'h20;
			14'd6937: ff_rdata <= 8'h01;
			14'd6938: ff_rdata <= 8'h0D;
			14'd6939: ff_rdata <= 8'h0D;
			14'd6940: ff_rdata <= 8'hC9;
			14'd6941: ff_rdata <= 8'hCD;
			14'd6942: ff_rdata <= 8'hF6;
			14'd6943: ff_rdata <= 8'h5A;
			14'd6944: ff_rdata <= 8'h2E;
			14'd6945: ff_rdata <= 8'h0F;
			14'd6946: ff_rdata <= 8'hCD;
			14'd6947: ff_rdata <= 8'hE4;
			14'd6948: ff_rdata <= 8'h67;
			14'd6949: ff_rdata <= 8'h5E;
			14'd6950: ff_rdata <= 8'h06;
			14'd6951: ff_rdata <= 8'h00;
			14'd6952: ff_rdata <= 8'h21;
			14'd6953: ff_rdata <= 8'h16;
			14'd6954: ff_rdata <= 8'h5A;
			14'd6955: ff_rdata <= 8'h09;
			14'd6956: ff_rdata <= 8'h4E;
			14'd6957: ff_rdata <= 8'h21;
			14'd6958: ff_rdata <= 8'h25;
			14'd6959: ff_rdata <= 8'h5A;
			14'd6960: ff_rdata <= 8'h09;
			14'd6961: ff_rdata <= 8'h7B;
			14'd6962: ff_rdata <= 8'h5E;
			14'd6963: ff_rdata <= 8'h23;
			14'd6964: ff_rdata <= 8'h56;
			14'd6965: ff_rdata <= 8'h3D;
			14'd6966: ff_rdata <= 8'h28;
			14'd6967: ff_rdata <= 8'h09;
			14'd6968: ff_rdata <= 8'hCB;
			14'd6969: ff_rdata <= 8'h3A;
			14'd6970: ff_rdata <= 8'hCB;
			14'd6971: ff_rdata <= 8'h1B;
			14'd6972: ff_rdata <= 8'h18;
			14'd6973: ff_rdata <= 8'hF7;
			14'd6974: ff_rdata <= 8'hCD;
			14'd6975: ff_rdata <= 8'h70;
			14'd6976: ff_rdata <= 8'h67;
			14'd6977: ff_rdata <= 8'h8B;
			14'd6978: ff_rdata <= 8'h5F;
			14'd6979: ff_rdata <= 8'h8A;
			14'd6980: ff_rdata <= 8'h93;
			14'd6981: ff_rdata <= 8'h57;
			14'd6982: ff_rdata <= 8'hD5;
			14'd6983: ff_rdata <= 8'h2E;
			14'd6984: ff_rdata <= 8'h10;
			14'd6985: ff_rdata <= 8'hCD;
			14'd6986: ff_rdata <= 8'hE4;
			14'd6987: ff_rdata <= 8'h67;
			14'd6988: ff_rdata <= 8'h4E;
			14'd6989: ff_rdata <= 8'hE5;
			14'd6990: ff_rdata <= 8'hCD;
			14'd6991: ff_rdata <= 8'h1A;
			14'd6992: ff_rdata <= 8'h66;
			14'd6993: ff_rdata <= 8'h28;
			14'd6994: ff_rdata <= 8'h11;
			14'd6995: ff_rdata <= 8'hC5;
			14'd6996: ff_rdata <= 8'hCD;
			14'd6997: ff_rdata <= 8'h51;
			14'd6998: ff_rdata <= 8'h66;
			14'd6999: ff_rdata <= 8'hC1;
			14'd7000: ff_rdata <= 8'h3E;
			14'd7001: ff_rdata <= 8'h40;
			14'd7002: ff_rdata <= 8'hBB;
			14'd7003: ff_rdata <= 8'h38;
			14'd7004: ff_rdata <= 8'hE1;
			14'd7005: ff_rdata <= 8'hCD;
			14'd7006: ff_rdata <= 8'h41;
			14'd7007: ff_rdata <= 8'h5C;
			14'd7008: ff_rdata <= 8'hB3;
			14'd7009: ff_rdata <= 8'h28;
			14'd7010: ff_rdata <= 8'h01;
			14'd7011: ff_rdata <= 8'h4B;
			14'd7012: ff_rdata <= 8'hE1;
			14'd7013: ff_rdata <= 8'h23;
			14'd7014: ff_rdata <= 8'hE5;
			14'd7015: ff_rdata <= 8'hCD;
			14'd7016: ff_rdata <= 8'hB0;
			14'd7017: ff_rdata <= 8'h5E;
			14'd7018: ff_rdata <= 8'hEB;
			14'd7019: ff_rdata <= 8'h01;
			14'd7020: ff_rdata <= 8'hF7;
			14'd7021: ff_rdata <= 8'hFF;
			14'd7022: ff_rdata <= 8'hE1;
			14'd7023: ff_rdata <= 8'hE5;
			14'd7024: ff_rdata <= 8'h09;
			14'd7025: ff_rdata <= 8'h72;
			14'd7026: ff_rdata <= 8'h23;
			14'd7027: ff_rdata <= 8'h73;
			14'd7028: ff_rdata <= 8'h23;
			14'd7029: ff_rdata <= 8'h0E;
			14'd7030: ff_rdata <= 8'h02;
			14'd7031: ff_rdata <= 8'hE3;
			14'd7032: ff_rdata <= 8'h23;
			14'd7033: ff_rdata <= 8'h5E;
			14'd7034: ff_rdata <= 8'h7B;
			14'd7035: ff_rdata <= 8'hE6;
			14'd7036: ff_rdata <= 8'hBF;
			14'd7037: ff_rdata <= 8'h77;
			14'd7038: ff_rdata <= 8'hE3;
			14'd7039: ff_rdata <= 8'h3E;
			14'd7040: ff_rdata <= 8'h80;
			14'd7041: ff_rdata <= 8'hB3;
			14'd7042: ff_rdata <= 8'h77;
			14'd7043: ff_rdata <= 8'h23;
			14'd7044: ff_rdata <= 8'h0C;
			14'd7045: ff_rdata <= 8'hE3;
			14'd7046: ff_rdata <= 8'h7B;
			14'd7047: ff_rdata <= 8'hE6;
			14'd7048: ff_rdata <= 8'h40;
			14'd7049: ff_rdata <= 8'h28;
			14'd7050: ff_rdata <= 8'h0C;
			14'd7051: ff_rdata <= 8'h23;
			14'd7052: ff_rdata <= 8'h5E;
			14'd7053: ff_rdata <= 8'h23;
			14'd7054: ff_rdata <= 8'h56;
			14'd7055: ff_rdata <= 8'hE1;
			14'd7056: ff_rdata <= 8'h72;
			14'd7057: ff_rdata <= 8'h23;
			14'd7058: ff_rdata <= 8'h73;
			14'd7059: ff_rdata <= 8'h23;
			14'd7060: ff_rdata <= 8'h0C;
			14'd7061: ff_rdata <= 8'h0C;
			14'd7062: ff_rdata <= 8'hFE;
			14'd7063: ff_rdata <= 8'hE1;
			14'd7064: ff_rdata <= 8'hD1;
			14'd7065: ff_rdata <= 8'h7A;
			14'd7066: ff_rdata <= 8'hB3;
			14'd7067: ff_rdata <= 8'h28;
			14'd7068: ff_rdata <= 8'h05;
			14'd7069: ff_rdata <= 8'h72;
			14'd7070: ff_rdata <= 8'h23;
			14'd7071: ff_rdata <= 8'h73;
			14'd7072: ff_rdata <= 8'h0C;
			14'd7073: ff_rdata <= 8'h0C;
			14'd7074: ff_rdata <= 8'h2E;
			14'd7075: ff_rdata <= 8'h07;
			14'd7076: ff_rdata <= 8'hCD;
			14'd7077: ff_rdata <= 8'hE4;
			14'd7078: ff_rdata <= 8'h67;
			14'd7079: ff_rdata <= 8'h71;
			14'd7080: ff_rdata <= 8'h79;
			14'd7081: ff_rdata <= 8'hD6;
			14'd7082: ff_rdata <= 8'h02;
			14'd7083: ff_rdata <= 8'h0F;
			14'd7084: ff_rdata <= 8'h0F;
			14'd7085: ff_rdata <= 8'h0F;
			14'd7086: ff_rdata <= 8'h23;
			14'd7087: ff_rdata <= 8'hB6;
			14'd7088: ff_rdata <= 8'h77;
			14'd7089: ff_rdata <= 8'h2B;
			14'd7090: ff_rdata <= 8'h7A;
			14'd7091: ff_rdata <= 8'hB3;
			14'd7092: ff_rdata <= 8'h20;
			14'd7093: ff_rdata <= 8'h0C;
			14'd7094: ff_rdata <= 8'hE5;
			14'd7095: ff_rdata <= 8'h3A;
			14'd7096: ff_rdata <= 8'h39;
			14'd7097: ff_rdata <= 8'hFB;
			14'd7098: ff_rdata <= 8'hF6;
			14'd7099: ff_rdata <= 8'h80;
			14'd7100: ff_rdata <= 8'h01;
			14'd7101: ff_rdata <= 8'h0B;
			14'd7102: ff_rdata <= 8'h00;
			14'd7103: ff_rdata <= 8'h09;
			14'd7104: ff_rdata <= 8'h77;
			14'd7105: ff_rdata <= 8'hE1;
			14'd7106: ff_rdata <= 8'hD1;
			14'd7107: ff_rdata <= 8'h46;
			14'd7108: ff_rdata <= 8'h23;
			14'd7109: ff_rdata <= 8'h5E;
			14'd7110: ff_rdata <= 8'h23;
			14'd7111: ff_rdata <= 8'hCD;
			14'd7112: ff_rdata <= 8'h9E;
			14'd7113: ff_rdata <= 8'h59;
			14'd7114: ff_rdata <= 8'h10;
			14'd7115: ff_rdata <= 8'hF9;
			14'd7116: ff_rdata <= 8'hCD;
			14'd7117: ff_rdata <= 8'hD5;
			14'd7118: ff_rdata <= 8'h59;
			14'd7119: ff_rdata <= 8'hDA;
			14'd7120: ff_rdata <= 8'h0F;
			14'd7121: ff_rdata <= 8'h59;
			14'd7122: ff_rdata <= 8'hC3;
			14'd7123: ff_rdata <= 8'hC6;
			14'd7124: ff_rdata <= 8'h65;
			14'd7125: ff_rdata <= 8'h44;
			14'd7126: ff_rdata <= 8'h4D;
			14'd7127: ff_rdata <= 8'hAF;
			14'd7128: ff_rdata <= 8'h67;
			14'd7129: ff_rdata <= 8'h6F;
			14'd7130: ff_rdata <= 8'hE5;
			14'd7131: ff_rdata <= 8'hED;
			14'd7132: ff_rdata <= 8'h42;
			14'd7133: ff_rdata <= 8'hEB;
			14'd7134: ff_rdata <= 8'h29;
			14'd7135: ff_rdata <= 8'h7C;
			14'd7136: ff_rdata <= 8'h4D;
			14'd7137: ff_rdata <= 8'hE1;
			14'd7138: ff_rdata <= 8'h06;
			14'd7139: ff_rdata <= 8'h10;
			14'd7140: ff_rdata <= 8'hED;
			14'd7141: ff_rdata <= 8'h6A;
			14'd7142: ff_rdata <= 8'h19;
			14'd7143: ff_rdata <= 8'h38;
			14'd7144: ff_rdata <= 8'h02;
			14'd7145: ff_rdata <= 8'hED;
			14'd7146: ff_rdata <= 8'h52;
			14'd7147: ff_rdata <= 8'hCB;
			14'd7148: ff_rdata <= 8'h11;
			14'd7149: ff_rdata <= 8'h17;
			14'd7150: ff_rdata <= 8'h10;
			14'd7151: ff_rdata <= 8'hF4;
			14'd7152: ff_rdata <= 8'h57;
			14'd7153: ff_rdata <= 8'h59;
			14'd7154: ff_rdata <= 8'hC9;
			14'd7155: ff_rdata <= 8'h1E;
			14'd7156: ff_rdata <= 8'h08;
			14'd7157: ff_rdata <= 8'h21;
			14'd7158: ff_rdata <= 8'h00;
			14'd7159: ff_rdata <= 8'h00;
			14'd7160: ff_rdata <= 8'h29;
			14'd7161: ff_rdata <= 8'h17;
			14'd7162: ff_rdata <= 8'h30;
			14'd7163: ff_rdata <= 8'h03;
			14'd7164: ff_rdata <= 8'h09;
			14'd7165: ff_rdata <= 8'hCE;
			14'd7166: ff_rdata <= 8'h00;
			14'd7167: ff_rdata <= 8'h1D;
			14'd7168: ff_rdata <= 8'hC2;
			14'd7169: ff_rdata <= 8'hF8;
			14'd7170: ff_rdata <= 8'h5B;
			14'd7171: ff_rdata <= 8'hC9;
			14'd7172: ff_rdata <= 8'h30;
			14'd7173: ff_rdata <= 8'h3E;
			14'd7174: ff_rdata <= 8'h7B;
			14'd7175: ff_rdata <= 8'hFE;
			14'd7176: ff_rdata <= 8'hC9;
			14'd7177: ff_rdata <= 8'h30;
			14'd7178: ff_rdata <= 8'h39;
			14'd7179: ff_rdata <= 8'hCD;
			14'd7180: ff_rdata <= 8'h41;
			14'd7181: ff_rdata <= 8'h5C;
			14'd7182: ff_rdata <= 8'hCD;
			14'd7183: ff_rdata <= 8'h1A;
			14'd7184: ff_rdata <= 8'h66;
			14'd7185: ff_rdata <= 8'hFE;
			14'd7186: ff_rdata <= 8'h2C;
			14'd7187: ff_rdata <= 8'h20;
			14'd7188: ff_rdata <= 8'h2F;
			14'd7189: ff_rdata <= 8'hCD;
			14'd7190: ff_rdata <= 8'h4E;
			14'd7191: ff_rdata <= 8'h66;
			14'd7192: ff_rdata <= 8'h18;
			14'd7193: ff_rdata <= 8'h27;
			14'd7194: ff_rdata <= 8'h38;
			14'd7195: ff_rdata <= 8'h02;
			14'd7196: ff_rdata <= 8'h1E;
			14'd7197: ff_rdata <= 8'h08;
			14'd7198: ff_rdata <= 8'h7B;
			14'd7199: ff_rdata <= 8'hFE;
			14'd7200: ff_rdata <= 8'h09;
			14'd7201: ff_rdata <= 8'h30;
			14'd7202: ff_rdata <= 8'h21;
			14'd7203: ff_rdata <= 8'h18;
			14'd7204: ff_rdata <= 8'h1C;
			14'd7205: ff_rdata <= 8'h30;
			14'd7206: ff_rdata <= 8'h1D;
			14'd7207: ff_rdata <= 8'h18;
			14'd7208: ff_rdata <= 8'h18;
			14'd7209: ff_rdata <= 8'hCD;
			14'd7210: ff_rdata <= 8'h14;
			14'd7211: ff_rdata <= 8'h66;
			14'd7212: ff_rdata <= 8'hFE;
			14'd7213: ff_rdata <= 8'h56;
			14'd7214: ff_rdata <= 8'h28;
			14'd7215: ff_rdata <= 8'h17;
			14'd7216: ff_rdata <= 8'hFE;
			14'd7217: ff_rdata <= 8'h57;
			14'd7218: ff_rdata <= 8'h28;
			14'd7219: ff_rdata <= 8'h26;
			14'd7220: ff_rdata <= 8'hCD;
			14'd7221: ff_rdata <= 8'h27;
			14'd7222: ff_rdata <= 8'h5D;
			14'd7223: ff_rdata <= 8'h38;
			14'd7224: ff_rdata <= 8'h0B;
			14'd7225: ff_rdata <= 8'hCD;
			14'd7226: ff_rdata <= 8'h51;
			14'd7227: ff_rdata <= 8'h66;
			14'd7228: ff_rdata <= 8'h7B;
			14'd7229: ff_rdata <= 8'hFE;
			14'd7230: ff_rdata <= 8'h40;
			14'd7231: ff_rdata <= 8'h30;
			14'd7232: ff_rdata <= 8'h03;
			14'd7233: ff_rdata <= 8'h7A;
			14'd7234: ff_rdata <= 8'hB7;
			14'd7235: ff_rdata <= 8'hC8;
			14'd7236: ff_rdata <= 8'hC3;
			14'd7237: ff_rdata <= 8'h70;
			14'd7238: ff_rdata <= 8'h67;
			14'd7239: ff_rdata <= 8'hCD;
			14'd7240: ff_rdata <= 8'h1A;
			14'd7241: ff_rdata <= 8'h66;
			14'd7242: ff_rdata <= 8'hC8;
			14'd7243: ff_rdata <= 8'hCD;
			14'd7244: ff_rdata <= 8'h27;
			14'd7245: ff_rdata <= 8'h5D;
			14'd7246: ff_rdata <= 8'h38;
			14'd7247: ff_rdata <= 8'hF4;
			14'd7248: ff_rdata <= 8'hCD;
			14'd7249: ff_rdata <= 8'h51;
			14'd7250: ff_rdata <= 8'h66;
			14'd7251: ff_rdata <= 8'h7B;
			14'd7252: ff_rdata <= 8'hFE;
			14'd7253: ff_rdata <= 8'h80;
			14'd7254: ff_rdata <= 8'h30;
			14'd7255: ff_rdata <= 8'hEC;
			14'd7256: ff_rdata <= 8'h18;
			14'd7257: ff_rdata <= 8'hE7;
			14'd7258: ff_rdata <= 8'hCD;
			14'd7259: ff_rdata <= 8'h1A;
			14'd7260: ff_rdata <= 8'h66;
			14'd7261: ff_rdata <= 8'h28;
			14'd7262: ff_rdata <= 8'h0E;
			14'd7263: ff_rdata <= 8'hCD;
			14'd7264: ff_rdata <= 8'h27;
			14'd7265: ff_rdata <= 8'h5D;
			14'd7266: ff_rdata <= 8'h38;
			14'd7267: ff_rdata <= 8'h06;
			14'd7268: ff_rdata <= 8'hCD;
			14'd7269: ff_rdata <= 8'h51;
			14'd7270: ff_rdata <= 8'h66;
			14'd7271: ff_rdata <= 8'hC3;
			14'd7272: ff_rdata <= 8'hB9;
			14'd7273: ff_rdata <= 8'h5A;
			14'd7274: ff_rdata <= 8'hCD;
			14'd7275: ff_rdata <= 8'h40;
			14'd7276: ff_rdata <= 8'h66;
			14'd7277: ff_rdata <= 8'hC3;
			14'd7278: ff_rdata <= 8'hB3;
			14'd7279: ff_rdata <= 8'h5A;
			14'd7280: ff_rdata <= 8'h41;
			14'd7281: ff_rdata <= 8'hED;
			14'd7282: ff_rdata <= 8'h5D;
			14'd7283: ff_rdata <= 8'h26;
			14'd7284: ff_rdata <= 8'h11;
			14'd7285: ff_rdata <= 8'h5F;
			14'd7286: ff_rdata <= 8'h7B;
			14'd7287: ff_rdata <= 8'h1A;
			14'd7288: ff_rdata <= 8'h5F;
			14'd7289: ff_rdata <= 8'hFD;
			14'd7290: ff_rdata <= 8'h96;
			14'd7291: ff_rdata <= 8'h5F;
			14'd7292: ff_rdata <= 8'hD9;
			14'd7293: ff_rdata <= 8'h37;
			14'd7294: ff_rdata <= 8'h5D;
			14'd7295: ff_rdata <= 8'hCC;
			14'd7296: ff_rdata <= 8'h80;
			14'd7297: ff_rdata <= 8'h5A;
			14'd7298: ff_rdata <= 8'hD1;
			14'd7299: ff_rdata <= 8'h9D;
			14'd7300: ff_rdata <= 8'h5D;
			14'd7301: ff_rdata <= 8'hD6;
			14'd7302: ff_rdata <= 8'h64;
			14'd7303: ff_rdata <= 8'h5D;
			14'd7304: ff_rdata <= 8'hCF;
			14'd7305: ff_rdata <= 8'hA6;
			14'd7306: ff_rdata <= 8'h5A;
			14'd7307: ff_rdata <= 8'h3E;
			14'd7308: ff_rdata <= 8'hAB;
			14'd7309: ff_rdata <= 8'h5D;
			14'd7310: ff_rdata <= 8'h3C;
			14'd7311: ff_rdata <= 8'hB8;
			14'd7312: ff_rdata <= 8'h5D;
			14'd7313: ff_rdata <= 8'hDA;
			14'd7314: ff_rdata <= 8'h61;
			14'd7315: ff_rdata <= 8'h5D;
			14'd7316: ff_rdata <= 8'h58;
			14'd7317: ff_rdata <= 8'hDB;
			14'd7318: ff_rdata <= 8'h66;
			14'd7319: ff_rdata <= 8'hD2;
			14'd7320: ff_rdata <= 8'hC3;
			14'd7321: ff_rdata <= 8'h5D;
			14'd7322: ff_rdata <= 8'hCE;
			14'd7323: ff_rdata <= 8'hE0;
			14'd7324: ff_rdata <= 8'h5D;
			14'd7325: ff_rdata <= 8'hD4;
			14'd7326: ff_rdata <= 8'h99;
			14'd7327: ff_rdata <= 8'h5A;
			14'd7328: ff_rdata <= 8'h40;
			14'd7329: ff_rdata <= 8'hAA;
			14'd7330: ff_rdata <= 8'h5C;
			14'd7331: ff_rdata <= 8'hCD;
			14'd7332: ff_rdata <= 8'h8E;
			14'd7333: ff_rdata <= 8'h5D;
			14'd7334: ff_rdata <= 8'hD3;
			14'd7335: ff_rdata <= 8'h95;
			14'd7336: ff_rdata <= 8'h5D;
			14'd7337: ff_rdata <= 8'h00;
			14'd7338: ff_rdata <= 8'hCD;
			14'd7339: ff_rdata <= 8'h14;
			14'd7340: ff_rdata <= 8'h66;
			14'd7341: ff_rdata <= 8'hFE;
			14'd7342: ff_rdata <= 8'h56;
			14'd7343: ff_rdata <= 8'h28;
			14'd7344: ff_rdata <= 8'h2C;
			14'd7345: ff_rdata <= 8'hFE;
			14'd7346: ff_rdata <= 8'h57;
			14'd7347: ff_rdata <= 8'h28;
			14'd7348: ff_rdata <= 8'h48;
			14'd7349: ff_rdata <= 8'hCD;
			14'd7350: ff_rdata <= 8'h27;
			14'd7351: ff_rdata <= 8'h5D;
			14'd7352: ff_rdata <= 8'h38;
			14'd7353: ff_rdata <= 8'h4C;
			14'd7354: ff_rdata <= 8'hCD;
			14'd7355: ff_rdata <= 8'h51;
			14'd7356: ff_rdata <= 8'h66;
			14'd7357: ff_rdata <= 8'hCD;
			14'd7358: ff_rdata <= 8'h41;
			14'd7359: ff_rdata <= 8'h5C;
			14'd7360: ff_rdata <= 8'h7B;
			14'd7361: ff_rdata <= 8'hFE;
			14'd7362: ff_rdata <= 8'h40;
			14'd7363: ff_rdata <= 8'h30;
			14'd7364: ff_rdata <= 8'h41;
			14'd7365: ff_rdata <= 8'h4F;
			14'd7366: ff_rdata <= 8'h3A;
			14'd7367: ff_rdata <= 8'h38;
			14'd7368: ff_rdata <= 8'hFB;
			14'd7369: ff_rdata <= 8'hCD;
			14'd7370: ff_rdata <= 8'h9F;
			14'd7371: ff_rdata <= 8'h61;
			14'd7372: ff_rdata <= 8'h30;
			14'd7373: ff_rdata <= 8'h05;
			14'd7374: ff_rdata <= 8'h79;
			14'd7375: ff_rdata <= 8'hFE;
			14'd7376: ff_rdata <= 8'h10;
			14'd7377: ff_rdata <= 8'h30;
			14'd7378: ff_rdata <= 8'h33;
			14'd7379: ff_rdata <= 8'h1E;
			14'd7380: ff_rdata <= 8'h84;
			14'd7381: ff_rdata <= 8'hCD;
			14'd7382: ff_rdata <= 8'hC5;
			14'd7383: ff_rdata <= 8'h59;
			14'd7384: ff_rdata <= 8'h59;
			14'd7385: ff_rdata <= 8'hC1;
			14'd7386: ff_rdata <= 8'hC3;
			14'd7387: ff_rdata <= 8'h75;
			14'd7388: ff_rdata <= 8'h5E;
			14'd7389: ff_rdata <= 8'hCD;
			14'd7390: ff_rdata <= 8'h14;
			14'd7391: ff_rdata <= 8'h66;
			14'd7392: ff_rdata <= 8'hCD;
			14'd7393: ff_rdata <= 8'h27;
			14'd7394: ff_rdata <= 8'h5D;
			14'd7395: ff_rdata <= 8'h38;
			14'd7396: ff_rdata <= 8'h21;
			14'd7397: ff_rdata <= 8'hCD;
			14'd7398: ff_rdata <= 8'h51;
			14'd7399: ff_rdata <= 8'h66;
			14'd7400: ff_rdata <= 8'h3E;
			14'd7401: ff_rdata <= 8'h7F;
			14'd7402: ff_rdata <= 8'h93;
			14'd7403: ff_rdata <= 8'hFA;
			14'd7404: ff_rdata <= 8'h06;
			14'd7405: ff_rdata <= 8'h5D;
			14'd7406: ff_rdata <= 8'h1F;
			14'd7407: ff_rdata <= 8'h4F;
			14'd7408: ff_rdata <= 8'hCD;
			14'd7409: ff_rdata <= 8'h41;
			14'd7410: ff_rdata <= 8'h5C;
			14'd7411: ff_rdata <= 8'h1E;
			14'd7412: ff_rdata <= 8'h85;
			14'd7413: ff_rdata <= 8'hCD;
			14'd7414: ff_rdata <= 8'hC5;
			14'd7415: ff_rdata <= 8'h59;
			14'd7416: ff_rdata <= 8'h59;
			14'd7417: ff_rdata <= 8'hC1;
			14'd7418: ff_rdata <= 8'hC3;
			14'd7419: ff_rdata <= 8'h75;
			14'd7420: ff_rdata <= 8'h5E;
			14'd7421: ff_rdata <= 8'hD1;
			14'd7422: ff_rdata <= 8'hCD;
			14'd7423: ff_rdata <= 8'h09;
			14'd7424: ff_rdata <= 8'h5D;
			14'd7425: ff_rdata <= 8'h1E;
			14'd7426: ff_rdata <= 8'h83;
			14'd7427: ff_rdata <= 8'hC3;
			14'd7428: ff_rdata <= 8'h6D;
			14'd7429: ff_rdata <= 8'h5E;
			14'd7430: ff_rdata <= 8'hC3;
			14'd7431: ff_rdata <= 8'h70;
			14'd7432: ff_rdata <= 8'h67;
			14'd7433: ff_rdata <= 8'hCD;
			14'd7434: ff_rdata <= 8'h82;
			14'd7435: ff_rdata <= 8'h5E;
			14'd7436: ff_rdata <= 8'hE5;
			14'd7437: ff_rdata <= 8'hCD;
			14'd7438: ff_rdata <= 8'h1A;
			14'd7439: ff_rdata <= 8'h66;
			14'd7440: ff_rdata <= 8'h28;
			14'd7441: ff_rdata <= 8'h11;
			14'd7442: ff_rdata <= 8'hC5;
			14'd7443: ff_rdata <= 8'hCD;
			14'd7444: ff_rdata <= 8'h51;
			14'd7445: ff_rdata <= 8'h66;
			14'd7446: ff_rdata <= 8'hC1;
			14'd7447: ff_rdata <= 8'h3E;
			14'd7448: ff_rdata <= 8'h40;
			14'd7449: ff_rdata <= 8'hBB;
			14'd7450: ff_rdata <= 8'h38;
			14'd7451: ff_rdata <= 8'hEA;
			14'd7452: ff_rdata <= 8'hCD;
			14'd7453: ff_rdata <= 8'h41;
			14'd7454: ff_rdata <= 8'h5C;
			14'd7455: ff_rdata <= 8'hB3;
			14'd7456: ff_rdata <= 8'h28;
			14'd7457: ff_rdata <= 8'hE4;
			14'd7458: ff_rdata <= 8'h4B;
			14'd7459: ff_rdata <= 8'hE1;
			14'd7460: ff_rdata <= 8'hC3;
			14'd7461: ff_rdata <= 8'hAF;
			14'd7462: ff_rdata <= 8'h5E;
			14'd7463: ff_rdata <= 8'hFE;
			14'd7464: ff_rdata <= 8'h2B;
			14'd7465: ff_rdata <= 8'hC8;
			14'd7466: ff_rdata <= 8'hFE;
			14'd7467: ff_rdata <= 8'h2D;
			14'd7468: ff_rdata <= 8'hC8;
			14'd7469: ff_rdata <= 8'hFE;
			14'd7470: ff_rdata <= 8'h3D;
			14'd7471: ff_rdata <= 8'hC8;
			14'd7472: ff_rdata <= 8'hFE;
			14'd7473: ff_rdata <= 8'h30;
			14'd7474: ff_rdata <= 8'hD8;
			14'd7475: ff_rdata <= 8'hFE;
			14'd7476: ff_rdata <= 8'h3A;
			14'd7477: ff_rdata <= 8'h3F;
			14'd7478: ff_rdata <= 8'hC9;
			14'd7479: ff_rdata <= 8'h30;
			14'd7480: ff_rdata <= 8'h28;
			14'd7481: ff_rdata <= 8'h7B;
			14'd7482: ff_rdata <= 8'hCD;
			14'd7483: ff_rdata <= 8'hF3;
			14'd7484: ff_rdata <= 8'h6D;
			14'd7485: ff_rdata <= 8'h38;
			14'd7486: ff_rdata <= 8'h22;
			14'd7487: ff_rdata <= 8'hCD;
			14'd7488: ff_rdata <= 8'h41;
			14'd7489: ff_rdata <= 8'h5C;
			14'd7490: ff_rdata <= 8'hD5;
			14'd7491: ff_rdata <= 8'hCD;
			14'd7492: ff_rdata <= 8'h14;
			14'd7493: ff_rdata <= 8'h66;
			14'd7494: ff_rdata <= 8'hFE;
			14'd7495: ff_rdata <= 8'h2C;
			14'd7496: ff_rdata <= 8'h20;
			14'd7497: ff_rdata <= 8'h17;
			14'd7498: ff_rdata <= 8'hCD;
			14'd7499: ff_rdata <= 8'h4E;
			14'd7500: ff_rdata <= 8'h66;
			14'd7501: ff_rdata <= 8'hCD;
			14'd7502: ff_rdata <= 8'h41;
			14'd7503: ff_rdata <= 8'h5C;
			14'd7504: ff_rdata <= 8'hD5;
			14'd7505: ff_rdata <= 8'h1E;
			14'd7506: ff_rdata <= 8'h82;
			14'd7507: ff_rdata <= 8'hCD;
			14'd7508: ff_rdata <= 8'hC5;
			14'd7509: ff_rdata <= 8'h59;
			14'd7510: ff_rdata <= 8'hE1;
			14'd7511: ff_rdata <= 8'hE3;
			14'd7512: ff_rdata <= 8'h5D;
			14'd7513: ff_rdata <= 8'hCD;
			14'd7514: ff_rdata <= 8'hC5;
			14'd7515: ff_rdata <= 8'h59;
			14'd7516: ff_rdata <= 8'hD1;
			14'd7517: ff_rdata <= 8'hC1;
			14'd7518: ff_rdata <= 8'hC3;
			14'd7519: ff_rdata <= 8'h75;
			14'd7520: ff_rdata <= 8'h5E;
			14'd7521: ff_rdata <= 8'hC3;
			14'd7522: ff_rdata <= 8'h70;
			14'd7523: ff_rdata <= 8'h67;
			14'd7524: ff_rdata <= 8'h38;
			14'd7525: ff_rdata <= 8'h02;
			14'd7526: ff_rdata <= 8'h1E;
			14'd7527: ff_rdata <= 8'h08;
			14'd7528: ff_rdata <= 8'hCD;
			14'd7529: ff_rdata <= 8'h41;
			14'd7530: ff_rdata <= 8'h5C;
			14'd7531: ff_rdata <= 8'h7B;
			14'd7532: ff_rdata <= 8'hFE;
			14'd7533: ff_rdata <= 8'h10;
			14'd7534: ff_rdata <= 8'h30;
			14'd7535: ff_rdata <= 8'h22;
			14'd7536: ff_rdata <= 8'h4F;
			14'd7537: ff_rdata <= 8'h1E;
			14'd7538: ff_rdata <= 8'h81;
			14'd7539: ff_rdata <= 8'hCD;
			14'd7540: ff_rdata <= 8'hC5;
			14'd7541: ff_rdata <= 8'h59;
			14'd7542: ff_rdata <= 8'h59;
			14'd7543: ff_rdata <= 8'hC1;
			14'd7544: ff_rdata <= 8'hC3;
			14'd7545: ff_rdata <= 8'h75;
			14'd7546: ff_rdata <= 8'h5E;
			14'd7547: ff_rdata <= 8'h38;
			14'd7548: ff_rdata <= 8'h02;
			14'd7549: ff_rdata <= 8'h1E;
			14'd7550: ff_rdata <= 8'h08;
			14'd7551: ff_rdata <= 8'hCD;
			14'd7552: ff_rdata <= 8'h41;
			14'd7553: ff_rdata <= 8'h5C;
			14'd7554: ff_rdata <= 8'h7B;
			14'd7555: ff_rdata <= 8'hFE;
			14'd7556: ff_rdata <= 8'h10;
			14'd7557: ff_rdata <= 8'h30;
			14'd7558: ff_rdata <= 8'h0B;
			14'd7559: ff_rdata <= 8'h3E;
			14'd7560: ff_rdata <= 8'h0F;
			14'd7561: ff_rdata <= 8'h93;
			14'd7562: ff_rdata <= 8'h87;
			14'd7563: ff_rdata <= 8'h5F;
			14'd7564: ff_rdata <= 8'h18;
			14'd7565: ff_rdata <= 8'hE2;
			14'd7566: ff_rdata <= 8'hD0;
			14'd7567: ff_rdata <= 8'h7B;
			14'd7568: ff_rdata <= 8'hB2;
			14'd7569: ff_rdata <= 8'hC0;
			14'd7570: ff_rdata <= 8'hC3;
			14'd7571: ff_rdata <= 8'h70;
			14'd7572: ff_rdata <= 8'h67;
			14'd7573: ff_rdata <= 8'h7B;
			14'd7574: ff_rdata <= 8'hFE;
			14'd7575: ff_rdata <= 8'h10;
			14'd7576: ff_rdata <= 8'h30;
			14'd7577: ff_rdata <= 8'hF8;
			14'd7578: ff_rdata <= 8'hC3;
			14'd7579: ff_rdata <= 8'h41;
			14'd7580: ff_rdata <= 8'h5C;
			14'd7581: ff_rdata <= 8'h38;
			14'd7582: ff_rdata <= 8'h02;
			14'd7583: ff_rdata <= 8'h1E;
			14'd7584: ff_rdata <= 8'h08;
			14'd7585: ff_rdata <= 8'h7B;
			14'd7586: ff_rdata <= 8'hFE;
			14'd7587: ff_rdata <= 8'h09;
			14'd7588: ff_rdata <= 8'h30;
			14'd7589: ff_rdata <= 8'hEC;
			14'd7590: ff_rdata <= 8'h2E;
			14'd7591: ff_rdata <= 8'h26;
			14'd7592: ff_rdata <= 8'hC3;
			14'd7593: ff_rdata <= 8'h8B;
			14'd7594: ff_rdata <= 8'h5A;
			14'd7595: ff_rdata <= 8'h2E;
			14'd7596: ff_rdata <= 8'h0F;
			14'd7597: ff_rdata <= 8'hCD;
			14'd7598: ff_rdata <= 8'hE4;
			14'd7599: ff_rdata <= 8'h67;
			14'd7600: ff_rdata <= 8'h7E;
			14'd7601: ff_rdata <= 8'h3C;
			14'd7602: ff_rdata <= 8'hFE;
			14'd7603: ff_rdata <= 8'h09;
			14'd7604: ff_rdata <= 8'h30;
			14'd7605: ff_rdata <= 8'hDC;
			14'd7606: ff_rdata <= 8'h77;
			14'd7607: ff_rdata <= 8'hC9;
			14'd7608: ff_rdata <= 8'h2E;
			14'd7609: ff_rdata <= 8'h0F;
			14'd7610: ff_rdata <= 8'hCD;
			14'd7611: ff_rdata <= 8'hE4;
			14'd7612: ff_rdata <= 8'h67;
			14'd7613: ff_rdata <= 8'h7E;
			14'd7614: ff_rdata <= 8'h3D;
			14'd7615: ff_rdata <= 8'h28;
			14'd7616: ff_rdata <= 8'hD1;
			14'd7617: ff_rdata <= 8'h77;
			14'd7618: ff_rdata <= 8'hC9;
			14'd7619: ff_rdata <= 8'h38;
			14'd7620: ff_rdata <= 8'h02;
			14'd7621: ff_rdata <= 8'h1E;
			14'd7622: ff_rdata <= 8'h04;
			14'd7623: ff_rdata <= 8'hCD;
			14'd7624: ff_rdata <= 8'h41;
			14'd7625: ff_rdata <= 8'h5C;
			14'd7626: ff_rdata <= 8'hB3;
			14'd7627: ff_rdata <= 8'h28;
			14'd7628: ff_rdata <= 8'hC5;
			14'd7629: ff_rdata <= 8'hFE;
			14'd7630: ff_rdata <= 8'h41;
			14'd7631: ff_rdata <= 8'h30;
			14'd7632: ff_rdata <= 8'hC1;
			14'd7633: ff_rdata <= 8'hAF;
			14'd7634: ff_rdata <= 8'hF5;
			14'd7635: ff_rdata <= 8'h21;
			14'd7636: ff_rdata <= 8'h11;
			14'd7637: ff_rdata <= 8'h5E;
			14'd7638: ff_rdata <= 8'hE5;
			14'd7639: ff_rdata <= 8'h2E;
			14'd7640: ff_rdata <= 8'h10;
			14'd7641: ff_rdata <= 8'hCD;
			14'd7642: ff_rdata <= 8'hE4;
			14'd7643: ff_rdata <= 8'h67;
			14'd7644: ff_rdata <= 8'hE5;
			14'd7645: ff_rdata <= 8'hC3;
			14'd7646: ff_rdata <= 8'hA2;
			14'd7647: ff_rdata <= 8'h5E;
			14'd7648: ff_rdata <= 8'h30;
			14'd7649: ff_rdata <= 8'hB0;
			14'd7650: ff_rdata <= 8'hCD;
			14'd7651: ff_rdata <= 8'h41;
			14'd7652: ff_rdata <= 8'h5C;
			14'd7653: ff_rdata <= 8'h7B;
			14'd7654: ff_rdata <= 8'hFE;
			14'd7655: ff_rdata <= 8'h61;
			14'd7656: ff_rdata <= 8'h38;
			14'd7657: ff_rdata <= 8'h1D;
			14'd7658: ff_rdata <= 8'hC3;
			14'd7659: ff_rdata <= 8'h70;
			14'd7660: ff_rdata <= 8'h67;
			14'd7661: ff_rdata <= 8'hCD;
			14'd7662: ff_rdata <= 8'hF6;
			14'd7663: ff_rdata <= 8'h5A;
			14'd7664: ff_rdata <= 8'h2E;
			14'd7665: ff_rdata <= 8'h0F;
			14'd7666: ff_rdata <= 8'hCD;
			14'd7667: ff_rdata <= 8'hE4;
			14'd7668: ff_rdata <= 8'h67;
			14'd7669: ff_rdata <= 8'h16;
			14'd7670: ff_rdata <= 8'h0C;
			14'd7671: ff_rdata <= 8'h46;
			14'd7672: ff_rdata <= 8'h3E;
			14'd7673: ff_rdata <= 8'hF4;
			14'd7674: ff_rdata <= 8'h82;
			14'd7675: ff_rdata <= 8'h10;
			14'd7676: ff_rdata <= 8'hFD;
			14'd7677: ff_rdata <= 8'h57;
			14'd7678: ff_rdata <= 8'h06;
			14'd7679: ff_rdata <= 8'h00;
			14'd7680: ff_rdata <= 8'h21;
			14'd7681: ff_rdata <= 8'h16;
			14'd7682: ff_rdata <= 8'h5A;
			14'd7683: ff_rdata <= 8'h09;
			14'd7684: ff_rdata <= 8'h7E;
			14'd7685: ff_rdata <= 8'h0F;
			14'd7686: ff_rdata <= 8'h82;
			14'd7687: ff_rdata <= 8'hC6;
			14'd7688: ff_rdata <= 8'h0C;
			14'd7689: ff_rdata <= 8'h57;
			14'd7690: ff_rdata <= 8'hCD;
			14'd7691: ff_rdata <= 8'h82;
			14'd7692: ff_rdata <= 8'h6C;
			14'd7693: ff_rdata <= 8'hD5;
			14'd7694: ff_rdata <= 8'hCD;
			14'd7695: ff_rdata <= 8'h94;
			14'd7696: ff_rdata <= 8'h5E;
			14'd7697: ff_rdata <= 8'hE5;
			14'd7698: ff_rdata <= 8'hCD;
			14'd7699: ff_rdata <= 8'h1A;
			14'd7700: ff_rdata <= 8'h66;
			14'd7701: ff_rdata <= 8'h28;
			14'd7702: ff_rdata <= 8'h09;
			14'd7703: ff_rdata <= 8'hFE;
			14'd7704: ff_rdata <= 8'h26;
			14'd7705: ff_rdata <= 8'hF5;
			14'd7706: ff_rdata <= 8'hCD;
			14'd7707: ff_rdata <= 8'h40;
			14'd7708: ff_rdata <= 8'h66;
			14'd7709: ff_rdata <= 8'hF1;
			14'd7710: ff_rdata <= 8'h28;
			14'd7711: ff_rdata <= 8'h41;
			14'd7712: ff_rdata <= 8'h2E;
			14'd7713: ff_rdata <= 8'h26;
			14'd7714: ff_rdata <= 8'hCD;
			14'd7715: ff_rdata <= 8'hE4;
			14'd7716: ff_rdata <= 8'h67;
			14'd7717: ff_rdata <= 8'h7E;
			14'd7718: ff_rdata <= 8'hFE;
			14'd7719: ff_rdata <= 8'h08;
			14'd7720: ff_rdata <= 8'h28;
			14'd7721: ff_rdata <= 8'h37;
			14'd7722: ff_rdata <= 8'hD1;
			14'd7723: ff_rdata <= 8'hD5;
			14'd7724: ff_rdata <= 8'h47;
			14'd7725: ff_rdata <= 8'h21;
			14'd7726: ff_rdata <= 8'h00;
			14'd7727: ff_rdata <= 8'h00;
			14'd7728: ff_rdata <= 8'h19;
			14'd7729: ff_rdata <= 8'h10;
			14'd7730: ff_rdata <= 8'hFD;
			14'd7731: ff_rdata <= 8'hCB;
			14'd7732: ff_rdata <= 8'h3C;
			14'd7733: ff_rdata <= 8'hCB;
			14'd7734: ff_rdata <= 8'h1D;
			14'd7735: ff_rdata <= 8'hCB;
			14'd7736: ff_rdata <= 8'h3C;
			14'd7737: ff_rdata <= 8'hCB;
			14'd7738: ff_rdata <= 8'h1D;
			14'd7739: ff_rdata <= 8'hCB;
			14'd7740: ff_rdata <= 8'h3C;
			14'd7741: ff_rdata <= 8'hCB;
			14'd7742: ff_rdata <= 8'h1D;
			14'd7743: ff_rdata <= 8'hD1;
			14'd7744: ff_rdata <= 8'hEB;
			14'd7745: ff_rdata <= 8'hB7;
			14'd7746: ff_rdata <= 8'hED;
			14'd7747: ff_rdata <= 8'h52;
			14'd7748: ff_rdata <= 8'hEB;
			14'd7749: ff_rdata <= 8'h28;
			14'd7750: ff_rdata <= 8'h1B;
			14'd7751: ff_rdata <= 8'hC1;
			14'd7752: ff_rdata <= 8'hF1;
			14'd7753: ff_rdata <= 8'hD5;
			14'd7754: ff_rdata <= 8'h58;
			14'd7755: ff_rdata <= 8'hCD;
			14'd7756: ff_rdata <= 8'hC5;
			14'd7757: ff_rdata <= 8'h59;
			14'd7758: ff_rdata <= 8'h78;
			14'd7759: ff_rdata <= 8'hB7;
			14'd7760: ff_rdata <= 8'h59;
			14'd7761: ff_rdata <= 8'hC4;
			14'd7762: ff_rdata <= 8'hC5;
			14'd7763: ff_rdata <= 8'h59;
			14'd7764: ff_rdata <= 8'h5D;
			14'd7765: ff_rdata <= 8'hCD;
			14'd7766: ff_rdata <= 8'hC5;
			14'd7767: ff_rdata <= 8'h59;
			14'd7768: ff_rdata <= 8'h5C;
			14'd7769: ff_rdata <= 8'hCD;
			14'd7770: ff_rdata <= 8'hC5;
			14'd7771: ff_rdata <= 8'h59;
			14'd7772: ff_rdata <= 8'hE1;
			14'd7773: ff_rdata <= 8'h1E;
			14'd7774: ff_rdata <= 8'h00;
			14'd7775: ff_rdata <= 8'h18;
			14'd7776: ff_rdata <= 8'h0C;
			14'd7777: ff_rdata <= 8'hE1;
			14'd7778: ff_rdata <= 8'hC1;
			14'd7779: ff_rdata <= 8'hD1;
			14'd7780: ff_rdata <= 8'h58;
			14'd7781: ff_rdata <= 8'hCD;
			14'd7782: ff_rdata <= 8'hC5;
			14'd7783: ff_rdata <= 8'h59;
			14'd7784: ff_rdata <= 8'h78;
			14'd7785: ff_rdata <= 8'hB7;
			14'd7786: ff_rdata <= 8'h28;
			14'd7787: ff_rdata <= 8'h04;
			14'd7788: ff_rdata <= 8'h59;
			14'd7789: ff_rdata <= 8'hCD;
			14'd7790: ff_rdata <= 8'hC5;
			14'd7791: ff_rdata <= 8'h59;
			14'd7792: ff_rdata <= 8'h5D;
			14'd7793: ff_rdata <= 8'hCD;
			14'd7794: ff_rdata <= 8'hC5;
			14'd7795: ff_rdata <= 8'h59;
			14'd7796: ff_rdata <= 8'h5C;
			14'd7797: ff_rdata <= 8'hCD;
			14'd7798: ff_rdata <= 8'hC5;
			14'd7799: ff_rdata <= 8'h59;
			14'd7800: ff_rdata <= 8'hCD;
			14'd7801: ff_rdata <= 8'hD5;
			14'd7802: ff_rdata <= 8'h59;
			14'd7803: ff_rdata <= 8'hFB;
			14'd7804: ff_rdata <= 8'hDA;
			14'd7805: ff_rdata <= 8'h0F;
			14'd7806: ff_rdata <= 8'h59;
			14'd7807: ff_rdata <= 8'hC3;
			14'd7808: ff_rdata <= 8'hC6;
			14'd7809: ff_rdata <= 8'h65;
			14'd7810: ff_rdata <= 8'h2E;
			14'd7811: ff_rdata <= 8'h09;
			14'd7812: ff_rdata <= 8'hCD;
			14'd7813: ff_rdata <= 8'hE4;
			14'd7814: ff_rdata <= 8'h67;
			14'd7815: ff_rdata <= 8'h4E;
			14'd7816: ff_rdata <= 8'h79;
			14'd7817: ff_rdata <= 8'hB7;
			14'd7818: ff_rdata <= 8'hF5;
			14'd7819: ff_rdata <= 8'h2E;
			14'd7820: ff_rdata <= 8'h10;
			14'd7821: ff_rdata <= 8'hCD;
			14'd7822: ff_rdata <= 8'hE4;
			14'd7823: ff_rdata <= 8'h67;
			14'd7824: ff_rdata <= 8'hF1;
			14'd7825: ff_rdata <= 8'hC0;
			14'd7826: ff_rdata <= 8'h4E;
			14'd7827: ff_rdata <= 8'hC9;
			14'd7828: ff_rdata <= 8'hCD;
			14'd7829: ff_rdata <= 8'h82;
			14'd7830: ff_rdata <= 8'h5E;
			14'd7831: ff_rdata <= 8'hE5;
			14'd7832: ff_rdata <= 8'hCD;
			14'd7833: ff_rdata <= 8'h1A;
			14'd7834: ff_rdata <= 8'h66;
			14'd7835: ff_rdata <= 8'h28;
			14'd7836: ff_rdata <= 8'h11;
			14'd7837: ff_rdata <= 8'hC5;
			14'd7838: ff_rdata <= 8'hCD;
			14'd7839: ff_rdata <= 8'h51;
			14'd7840: ff_rdata <= 8'h66;
			14'd7841: ff_rdata <= 8'hC1;
			14'd7842: ff_rdata <= 8'h3E;
			14'd7843: ff_rdata <= 8'h40;
			14'd7844: ff_rdata <= 8'hBB;
			14'd7845: ff_rdata <= 8'h38;
			14'd7846: ff_rdata <= 8'h70;
			14'd7847: ff_rdata <= 8'hCD;
			14'd7848: ff_rdata <= 8'h41;
			14'd7849: ff_rdata <= 8'h5C;
			14'd7850: ff_rdata <= 8'hB3;
			14'd7851: ff_rdata <= 8'h28;
			14'd7852: ff_rdata <= 8'h01;
			14'd7853: ff_rdata <= 8'h4B;
			14'd7854: ff_rdata <= 8'hE1;
			14'd7855: ff_rdata <= 8'h23;
			14'd7856: ff_rdata <= 8'h7E;
			14'd7857: ff_rdata <= 8'h06;
			14'd7858: ff_rdata <= 8'h00;
			14'd7859: ff_rdata <= 8'hCD;
			14'd7860: ff_rdata <= 8'hF3;
			14'd7861: ff_rdata <= 8'h5B;
			14'd7862: ff_rdata <= 8'hE5;
			14'd7863: ff_rdata <= 8'hED;
			14'd7864: ff_rdata <= 8'h5B;
			14'd7865: ff_rdata <= 8'h7A;
			14'd7866: ff_rdata <= 8'hF9;
			14'd7867: ff_rdata <= 8'hCD;
			14'd7868: ff_rdata <= 8'hD5;
			14'd7869: ff_rdata <= 8'h5B;
			14'd7870: ff_rdata <= 8'hEB;
			14'd7871: ff_rdata <= 8'hE3;
			14'd7872: ff_rdata <= 8'h06;
			14'd7873: ff_rdata <= 8'h05;
			14'd7874: ff_rdata <= 8'hCB;
			14'd7875: ff_rdata <= 8'h3C;
			14'd7876: ff_rdata <= 8'hCB;
			14'd7877: ff_rdata <= 8'h1D;
			14'd7878: ff_rdata <= 8'h10;
			14'd7879: ff_rdata <= 8'hFA;
			14'd7880: ff_rdata <= 8'hCD;
			14'd7881: ff_rdata <= 8'hD5;
			14'd7882: ff_rdata <= 8'h5B;
			14'd7883: ff_rdata <= 8'hCD;
			14'd7884: ff_rdata <= 8'h02;
			14'd7885: ff_rdata <= 8'h5F;
			14'd7886: ff_rdata <= 8'hDD;
			14'd7887: ff_rdata <= 8'h6E;
			14'd7888: ff_rdata <= 8'h00;
			14'd7889: ff_rdata <= 8'h26;
			14'd7890: ff_rdata <= 8'h00;
			14'd7891: ff_rdata <= 8'h19;
			14'd7892: ff_rdata <= 8'hDD;
			14'd7893: ff_rdata <= 8'h75;
			14'd7894: ff_rdata <= 8'h00;
			14'd7895: ff_rdata <= 8'h11;
			14'd7896: ff_rdata <= 8'hE0;
			14'd7897: ff_rdata <= 8'hFF;
			14'd7898: ff_rdata <= 8'h19;
			14'd7899: ff_rdata <= 8'h30;
			14'd7900: ff_rdata <= 8'h06;
			14'd7901: ff_rdata <= 8'hDD;
			14'd7902: ff_rdata <= 8'h75;
			14'd7903: ff_rdata <= 8'h00;
			14'd7904: ff_rdata <= 8'hE1;
			14'd7905: ff_rdata <= 8'h23;
			14'd7906: ff_rdata <= 8'hE5;
			14'd7907: ff_rdata <= 8'hD1;
			14'd7908: ff_rdata <= 8'h62;
			14'd7909: ff_rdata <= 8'h6B;
			14'd7910: ff_rdata <= 8'hCD;
			14'd7911: ff_rdata <= 8'h1A;
			14'd7912: ff_rdata <= 8'h66;
			14'd7913: ff_rdata <= 8'h28;
			14'd7914: ff_rdata <= 8'h16;
			14'd7915: ff_rdata <= 8'hFE;
			14'd7916: ff_rdata <= 8'h2E;
			14'd7917: ff_rdata <= 8'h20;
			14'd7918: ff_rdata <= 8'h0F;
			14'd7919: ff_rdata <= 8'hCB;
			14'd7920: ff_rdata <= 8'h3A;
			14'd7921: ff_rdata <= 8'hCB;
			14'd7922: ff_rdata <= 8'h1B;
			14'd7923: ff_rdata <= 8'hED;
			14'd7924: ff_rdata <= 8'h5A;
			14'd7925: ff_rdata <= 8'h3E;
			14'd7926: ff_rdata <= 8'hE0;
			14'd7927: ff_rdata <= 8'hA4;
			14'd7928: ff_rdata <= 8'h28;
			14'd7929: ff_rdata <= 8'hEC;
			14'd7930: ff_rdata <= 8'hAC;
			14'd7931: ff_rdata <= 8'h67;
			14'd7932: ff_rdata <= 8'h18;
			14'd7933: ff_rdata <= 8'h03;
			14'd7934: ff_rdata <= 8'hCD;
			14'd7935: ff_rdata <= 8'h40;
			14'd7936: ff_rdata <= 8'h66;
			14'd7937: ff_rdata <= 8'hC9;
			14'd7938: ff_rdata <= 8'hC5;
			14'd7939: ff_rdata <= 8'h3A;
			14'd7940: ff_rdata <= 8'h38;
			14'd7941: ff_rdata <= 8'hFB;
			14'd7942: ff_rdata <= 8'h4F;
			14'd7943: ff_rdata <= 8'h06;
			14'd7944: ff_rdata <= 8'h00;
			14'd7945: ff_rdata <= 8'hDD;
			14'd7946: ff_rdata <= 8'h21;
			14'd7947: ff_rdata <= 8'h19;
			14'd7948: ff_rdata <= 8'hFA;
			14'd7949: ff_rdata <= 8'hDD;
			14'd7950: ff_rdata <= 8'h09;
			14'd7951: ff_rdata <= 8'hC1;
			14'd7952: ff_rdata <= 8'hC9;
			14'd7953: ff_rdata <= 8'h1E;
			14'd7954: ff_rdata <= 8'h87;
			14'd7955: ff_rdata <= 8'hC1;
			14'd7956: ff_rdata <= 8'hC3;
			14'd7957: ff_rdata <= 8'h75;
			14'd7958: ff_rdata <= 8'h5E;
			14'd7959: ff_rdata <= 8'hC3;
			14'd7960: ff_rdata <= 8'h70;
			14'd7961: ff_rdata <= 8'h67;
			14'd7962: ff_rdata <= 8'h2E;
			14'd7963: ff_rdata <= 8'h09;
			14'd7964: ff_rdata <= 8'hCD;
			14'd7965: ff_rdata <= 8'hE4;
			14'd7966: ff_rdata <= 8'h67;
			14'd7967: ff_rdata <= 8'h7E;
			14'd7968: ff_rdata <= 8'h20;
			14'd7969: ff_rdata <= 8'hF5;
			14'd7970: ff_rdata <= 8'h0E;
			14'd7971: ff_rdata <= 8'h00;
			14'd7972: ff_rdata <= 8'h2A;
			14'd7973: ff_rdata <= 8'h3C;
			14'd7974: ff_rdata <= 8'hFB;
			14'd7975: ff_rdata <= 8'hE5;
			14'd7976: ff_rdata <= 8'h3A;
			14'd7977: ff_rdata <= 8'h3B;
			14'd7978: ff_rdata <= 8'hFB;
			14'd7979: ff_rdata <= 8'hF5;
			14'd7980: ff_rdata <= 8'hCD;
			14'd7981: ff_rdata <= 8'h14;
			14'd7982: ff_rdata <= 8'h66;
			14'd7983: ff_rdata <= 8'hFE;
			14'd7984: ff_rdata <= 8'h4E;
			14'd7985: ff_rdata <= 8'h28;
			14'd7986: ff_rdata <= 8'h0C;
			14'd7987: ff_rdata <= 8'hFE;
			14'd7988: ff_rdata <= 8'h52;
			14'd7989: ff_rdata <= 8'h28;
			14'd7990: ff_rdata <= 8'h08;
			14'd7991: ff_rdata <= 8'hFE;
			14'd7992: ff_rdata <= 8'h41;
			14'd7993: ff_rdata <= 8'h38;
			14'd7994: ff_rdata <= 8'h07;
			14'd7995: ff_rdata <= 8'hFE;
			14'd7996: ff_rdata <= 8'h48;
			14'd7997: ff_rdata <= 8'h30;
			14'd7998: ff_rdata <= 8'h03;
			14'd7999: ff_rdata <= 8'h0C;
			14'd8000: ff_rdata <= 8'h18;
			14'd8001: ff_rdata <= 8'hEA;
			14'd8002: ff_rdata <= 8'hFE;
			14'd8003: ff_rdata <= 8'h7D;
			14'd8004: ff_rdata <= 8'h28;
			14'd8005: ff_rdata <= 8'h0F;
			14'd8006: ff_rdata <= 8'hFE;
			14'd8007: ff_rdata <= 8'h7B;
			14'd8008: ff_rdata <= 8'h28;
			14'd8009: ff_rdata <= 8'hCD;
			14'd8010: ff_rdata <= 8'hFE;
			14'd8011: ff_rdata <= 8'h3D;
			14'd8012: ff_rdata <= 8'h20;
			14'd8013: ff_rdata <= 8'hDE;
			14'd8014: ff_rdata <= 8'hC5;
			14'd8015: ff_rdata <= 8'hCD;
			14'd8016: ff_rdata <= 8'hA4;
			14'd8017: ff_rdata <= 8'h66;
			14'd8018: ff_rdata <= 8'hC1;
			14'd8019: ff_rdata <= 8'h18;
			14'd8020: ff_rdata <= 8'hDA;
			14'd8021: ff_rdata <= 8'h2E;
			14'd8022: ff_rdata <= 8'h10;
			14'd8023: ff_rdata <= 8'hCD;
			14'd8024: ff_rdata <= 8'hE4;
			14'd8025: ff_rdata <= 8'h67;
			14'd8026: ff_rdata <= 8'h5E;
			14'd8027: ff_rdata <= 8'h16;
			14'd8028: ff_rdata <= 8'h00;
			14'd8029: ff_rdata <= 8'hCD;
			14'd8030: ff_rdata <= 8'h1A;
			14'd8031: ff_rdata <= 8'h66;
			14'd8032: ff_rdata <= 8'h28;
			14'd8033: ff_rdata <= 8'h0D;
			14'd8034: ff_rdata <= 8'hCD;
			14'd8035: ff_rdata <= 8'h40;
			14'd8036: ff_rdata <= 8'h66;
			14'd8037: ff_rdata <= 8'hCD;
			14'd8038: ff_rdata <= 8'h27;
			14'd8039: ff_rdata <= 8'h5D;
			14'd8040: ff_rdata <= 8'h38;
			14'd8041: ff_rdata <= 8'h05;
			14'd8042: ff_rdata <= 8'hC5;
			14'd8043: ff_rdata <= 8'hCD;
			14'd8044: ff_rdata <= 8'h4E;
			14'd8045: ff_rdata <= 8'h66;
			14'd8046: ff_rdata <= 8'hC1;
			14'd8047: ff_rdata <= 8'h3E;
			14'd8048: ff_rdata <= 8'h40;
			14'd8049: ff_rdata <= 8'hBB;
			14'd8050: ff_rdata <= 8'h38;
			14'd8051: ff_rdata <= 8'hA3;
			14'd8052: ff_rdata <= 8'hCD;
			14'd8053: ff_rdata <= 8'h41;
			14'd8054: ff_rdata <= 8'h5C;
			14'd8055: ff_rdata <= 8'h79;
			14'd8056: ff_rdata <= 8'h42;
			14'd8057: ff_rdata <= 8'h4B;
			14'd8058: ff_rdata <= 8'hCD;
			14'd8059: ff_rdata <= 8'hF3;
			14'd8060: ff_rdata <= 8'h5B;
			14'd8061: ff_rdata <= 8'hB4;
			14'd8062: ff_rdata <= 8'h20;
			14'd8063: ff_rdata <= 8'h97;
			14'd8064: ff_rdata <= 8'h7D;
			14'd8065: ff_rdata <= 8'hFE;
			14'd8066: ff_rdata <= 8'h41;
			14'd8067: ff_rdata <= 8'h30;
			14'd8068: ff_rdata <= 8'h92;
			14'd8069: ff_rdata <= 8'hF5;
			14'd8070: ff_rdata <= 8'h2E;
			14'd8071: ff_rdata <= 8'h09;
			14'd8072: ff_rdata <= 8'hCD;
			14'd8073: ff_rdata <= 8'hE4;
			14'd8074: ff_rdata <= 8'h67;
			14'd8075: ff_rdata <= 8'hF1;
			14'd8076: ff_rdata <= 8'h77;
			14'd8077: ff_rdata <= 8'hF1;
			14'd8078: ff_rdata <= 8'h32;
			14'd8079: ff_rdata <= 8'h3B;
			14'd8080: ff_rdata <= 8'hFB;
			14'd8081: ff_rdata <= 8'hE1;
			14'd8082: ff_rdata <= 8'h22;
			14'd8083: ff_rdata <= 8'h3C;
			14'd8084: ff_rdata <= 8'hFB;
			14'd8085: ff_rdata <= 8'hC9;
			14'd8086: ff_rdata <= 8'h2E;
			14'd8087: ff_rdata <= 8'h09;
			14'd8088: ff_rdata <= 8'hCD;
			14'd8089: ff_rdata <= 8'hE4;
			14'd8090: ff_rdata <= 8'h67;
			14'd8091: ff_rdata <= 8'h7E;
			14'd8092: ff_rdata <= 8'hB7;
			14'd8093: ff_rdata <= 8'h28;
			14'd8094: ff_rdata <= 8'h2F;
			14'd8095: ff_rdata <= 8'h36;
			14'd8096: ff_rdata <= 8'h00;
			14'd8097: ff_rdata <= 8'hC9;
			14'd8098: ff_rdata <= 8'h42;
			14'd8099: ff_rdata <= 8'hD1;
			14'd8100: ff_rdata <= 8'h5F;
			14'd8101: ff_rdata <= 8'h53;
			14'd8102: ff_rdata <= 8'hD1;
			14'd8103: ff_rdata <= 8'h5F;
			14'd8104: ff_rdata <= 8'h4D;
			14'd8105: ff_rdata <= 8'hD1;
			14'd8106: ff_rdata <= 8'h5F;
			14'd8107: ff_rdata <= 8'h43;
			14'd8108: ff_rdata <= 8'hD1;
			14'd8109: ff_rdata <= 8'h5F;
			14'd8110: ff_rdata <= 8'h48;
			14'd8111: ff_rdata <= 8'hD1;
			14'd8112: ff_rdata <= 8'h5F;
			14'd8113: ff_rdata <= 8'hD2;
			14'd8114: ff_rdata <= 8'hC3;
			14'd8115: ff_rdata <= 8'h5D;
			14'd8116: ff_rdata <= 8'h40;
			14'd8117: ff_rdata <= 8'h2A;
			14'd8118: ff_rdata <= 8'h60;
			14'd8119: ff_rdata <= 8'hD4;
			14'd8120: ff_rdata <= 8'h99;
			14'd8121: ff_rdata <= 8'h5A;
			14'd8122: ff_rdata <= 8'hD9;
			14'd8123: ff_rdata <= 8'h37;
			14'd8124: ff_rdata <= 8'h5D;
			14'd8125: ff_rdata <= 8'hD6;
			14'd8126: ff_rdata <= 8'h7B;
			14'd8127: ff_rdata <= 8'h5D;
			14'd8128: ff_rdata <= 8'h58;
			14'd8129: ff_rdata <= 8'hDB;
			14'd8130: ff_rdata <= 8'h66;
			14'd8131: ff_rdata <= 8'h00;
			14'd8132: ff_rdata <= 8'h42;
			14'd8133: ff_rdata <= 8'h53;
			14'd8134: ff_rdata <= 8'h4D;
			14'd8135: ff_rdata <= 8'h43;
			14'd8136: ff_rdata <= 8'h48;
			14'd8137: ff_rdata <= 8'h10;
			14'd8138: ff_rdata <= 8'h08;
			14'd8139: ff_rdata <= 8'h04;
			14'd8140: ff_rdata <= 8'h02;
			14'd8141: ff_rdata <= 8'h01;
			14'd8142: ff_rdata <= 8'hC3;
			14'd8143: ff_rdata <= 8'h70;
			14'd8144: ff_rdata <= 8'h67;
			14'd8145: ff_rdata <= 8'h01;
			14'd8146: ff_rdata <= 8'h00;
			14'd8147: ff_rdata <= 8'h00;
			14'd8148: ff_rdata <= 8'hCD;
			14'd8149: ff_rdata <= 8'h40;
			14'd8150: ff_rdata <= 8'h66;
			14'd8151: ff_rdata <= 8'hCD;
			14'd8152: ff_rdata <= 8'h14;
			14'd8153: ff_rdata <= 8'h66;
			14'd8154: ff_rdata <= 8'hCD;
			14'd8155: ff_rdata <= 8'h27;
			14'd8156: ff_rdata <= 8'h5D;
			14'd8157: ff_rdata <= 8'h30;
			14'd8158: ff_rdata <= 8'h24;
			14'd8159: ff_rdata <= 8'hC5;
			14'd8160: ff_rdata <= 8'h21;
			14'd8161: ff_rdata <= 8'hC4;
			14'd8162: ff_rdata <= 8'h5F;
			14'd8163: ff_rdata <= 8'h01;
			14'd8164: ff_rdata <= 8'h05;
			14'd8165: ff_rdata <= 8'h00;
			14'd8166: ff_rdata <= 8'hED;
			14'd8167: ff_rdata <= 8'hB1;
			14'd8168: ff_rdata <= 8'h20;
			14'd8169: ff_rdata <= 8'hE4;
			14'd8170: ff_rdata <= 8'h0E;
			14'd8171: ff_rdata <= 8'h04;
			14'd8172: ff_rdata <= 8'h09;
			14'd8173: ff_rdata <= 8'h56;
			14'd8174: ff_rdata <= 8'hC1;
			14'd8175: ff_rdata <= 8'hCD;
			14'd8176: ff_rdata <= 8'h14;
			14'd8177: ff_rdata <= 8'h66;
			14'd8178: ff_rdata <= 8'hFE;
			14'd8179: ff_rdata <= 8'h21;
			14'd8180: ff_rdata <= 8'hF5;
			14'd8181: ff_rdata <= 8'hC4;
			14'd8182: ff_rdata <= 8'h40;
			14'd8183: ff_rdata <= 8'h66;
			14'd8184: ff_rdata <= 8'hF1;
			14'd8185: ff_rdata <= 8'h20;
			14'd8186: ff_rdata <= 8'h03;
			14'd8187: ff_rdata <= 8'h7A;
			14'd8188: ff_rdata <= 8'hB0;
			14'd8189: ff_rdata <= 8'h47;
			14'd8190: ff_rdata <= 8'h7A;
			14'd8191: ff_rdata <= 8'hB1;
			14'd8192: ff_rdata <= 8'h4F;
			14'd8193: ff_rdata <= 8'h18;
			14'd8194: ff_rdata <= 8'hD4;
			14'd8195: ff_rdata <= 8'h0C;
			14'd8196: ff_rdata <= 8'h0D;
			14'd8197: ff_rdata <= 8'h28;
			14'd8198: ff_rdata <= 8'hC7;
			14'd8199: ff_rdata <= 8'h3E;
			14'd8200: ff_rdata <= 8'hC0;
			14'd8201: ff_rdata <= 8'hB1;
			14'd8202: ff_rdata <= 8'hF5;
			14'd8203: ff_rdata <= 8'hC5;
			14'd8204: ff_rdata <= 8'h21;
			14'd8205: ff_rdata <= 8'h1F;
			14'd8206: ff_rdata <= 8'h60;
			14'd8207: ff_rdata <= 8'hE5;
			14'd8208: ff_rdata <= 8'h2E;
			14'd8209: ff_rdata <= 8'h10;
			14'd8210: ff_rdata <= 8'hCD;
			14'd8211: ff_rdata <= 8'hE4;
			14'd8212: ff_rdata <= 8'h67;
			14'd8213: ff_rdata <= 8'hE5;
			14'd8214: ff_rdata <= 8'hCD;
			14'd8215: ff_rdata <= 8'h40;
			14'd8216: ff_rdata <= 8'h66;
			14'd8217: ff_rdata <= 8'hCD;
			14'd8218: ff_rdata <= 8'h4E;
			14'd8219: ff_rdata <= 8'h66;
			14'd8220: ff_rdata <= 8'hC3;
			14'd8221: ff_rdata <= 8'hA2;
			14'd8222: ff_rdata <= 8'h5E;
			14'd8223: ff_rdata <= 8'hC1;
			14'd8224: ff_rdata <= 8'hF1;
			14'd8225: ff_rdata <= 8'hD1;
			14'd8226: ff_rdata <= 8'h5F;
			14'd8227: ff_rdata <= 8'hCD;
			14'd8228: ff_rdata <= 8'hC5;
			14'd8229: ff_rdata <= 8'h59;
			14'd8230: ff_rdata <= 8'h58;
			14'd8231: ff_rdata <= 8'hC3;
			14'd8232: ff_rdata <= 8'h6D;
			14'd8233: ff_rdata <= 8'h5E;
			14'd8234: ff_rdata <= 8'hCD;
			14'd8235: ff_rdata <= 8'h14;
			14'd8236: ff_rdata <= 8'h66;
			14'd8237: ff_rdata <= 8'hFE;
			14'd8238: ff_rdata <= 8'h56;
			14'd8239: ff_rdata <= 8'hCA;
			14'd8240: ff_rdata <= 8'hDD;
			14'd8241: ff_rdata <= 8'h5C;
			14'd8242: ff_rdata <= 8'hFE;
			14'd8243: ff_rdata <= 8'h41;
			14'd8244: ff_rdata <= 8'h20;
			14'd8245: ff_rdata <= 8'h98;
			14'd8246: ff_rdata <= 8'hCD;
			14'd8247: ff_rdata <= 8'h14;
			14'd8248: ff_rdata <= 8'h66;
			14'd8249: ff_rdata <= 8'hCD;
			14'd8250: ff_rdata <= 8'h27;
			14'd8251: ff_rdata <= 8'h5D;
			14'd8252: ff_rdata <= 8'h38;
			14'd8253: ff_rdata <= 8'h1A;
			14'd8254: ff_rdata <= 8'hCD;
			14'd8255: ff_rdata <= 8'h51;
			14'd8256: ff_rdata <= 8'h66;
			14'd8257: ff_rdata <= 8'hCD;
			14'd8258: ff_rdata <= 8'h41;
			14'd8259: ff_rdata <= 8'h5C;
			14'd8260: ff_rdata <= 8'h7B;
			14'd8261: ff_rdata <= 8'hFE;
			14'd8262: ff_rdata <= 8'h10;
			14'd8263: ff_rdata <= 8'h30;
			14'd8264: ff_rdata <= 8'h0F;
			14'd8265: ff_rdata <= 8'h3E;
			14'd8266: ff_rdata <= 8'h0F;
			14'd8267: ff_rdata <= 8'h93;
			14'd8268: ff_rdata <= 8'h87;
			14'd8269: ff_rdata <= 8'h4F;
			14'd8270: ff_rdata <= 8'h1E;
			14'd8271: ff_rdata <= 8'h86;
			14'd8272: ff_rdata <= 8'hCD;
			14'd8273: ff_rdata <= 8'hC5;
			14'd8274: ff_rdata <= 8'h59;
			14'd8275: ff_rdata <= 8'h59;
			14'd8276: ff_rdata <= 8'hC1;
			14'd8277: ff_rdata <= 8'hC3;
			14'd8278: ff_rdata <= 8'h75;
			14'd8279: ff_rdata <= 8'h5E;
			14'd8280: ff_rdata <= 8'hC3;
			14'd8281: ff_rdata <= 8'h70;
			14'd8282: ff_rdata <= 8'h67;
			14'd8283: ff_rdata <= 8'hF5;
			14'd8284: ff_rdata <= 8'hF3;
			14'd8285: ff_rdata <= 8'h21;
			14'd8286: ff_rdata <= 8'h99;
			14'd8287: ff_rdata <= 8'hF9;
			14'd8288: ff_rdata <= 8'h3A;
			14'd8289: ff_rdata <= 8'h83;
			14'd8290: ff_rdata <= 8'hF9;
			14'd8291: ff_rdata <= 8'hB7;
			14'd8292: ff_rdata <= 8'h20;
			14'd8293: ff_rdata <= 8'h1C;
			14'd8294: ff_rdata <= 8'h2F;
			14'd8295: ff_rdata <= 8'h32;
			14'd8296: ff_rdata <= 8'h83;
			14'd8297: ff_rdata <= 8'hF9;
			14'd8298: ff_rdata <= 8'hE5;
			14'd8299: ff_rdata <= 8'hAF;
			14'd8300: ff_rdata <= 8'h32;
			14'd8301: ff_rdata <= 8'h26;
			14'd8302: ff_rdata <= 8'hFA;
			14'd8303: ff_rdata <= 8'hCD;
			14'd8304: ff_rdata <= 8'h87;
			14'd8305: ff_rdata <= 8'h60;
			14'd8306: ff_rdata <= 8'h3A;
			14'd8307: ff_rdata <= 8'h26;
			14'd8308: ff_rdata <= 8'hFA;
			14'd8309: ff_rdata <= 8'hB7;
			14'd8310: ff_rdata <= 8'h20;
			14'd8311: ff_rdata <= 8'hF3;
			14'd8312: ff_rdata <= 8'hE1;
			14'd8313: ff_rdata <= 8'hF3;
			14'd8314: ff_rdata <= 8'hAF;
			14'd8315: ff_rdata <= 8'h32;
			14'd8316: ff_rdata <= 8'h83;
			14'd8317: ff_rdata <= 8'hF9;
			14'd8318: ff_rdata <= 8'h35;
			14'd8319: ff_rdata <= 8'hF2;
			14'd8320: ff_rdata <= 8'h66;
			14'd8321: ff_rdata <= 8'h60;
			14'd8322: ff_rdata <= 8'h34;
			14'd8323: ff_rdata <= 8'hF1;
			14'd8324: ff_rdata <= 8'hC3;
			14'd8325: ff_rdata <= 8'hBB;
			14'd8326: ff_rdata <= 8'hF9;
			14'd8327: ff_rdata <= 8'h3A;
			14'd8328: ff_rdata <= 8'h3F;
			14'd8329: ff_rdata <= 8'hFB;
			14'd8330: ff_rdata <= 8'hB7;
			14'd8331: ff_rdata <= 8'h28;
			14'd8332: ff_rdata <= 8'h0A;
			14'd8333: ff_rdata <= 8'hCD;
			14'd8334: ff_rdata <= 8'hB1;
			14'd8335: ff_rdata <= 8'h63;
			14'd8336: ff_rdata <= 8'h20;
			14'd8337: ff_rdata <= 8'h12;
			14'd8338: ff_rdata <= 8'h3A;
			14'd8339: ff_rdata <= 8'h3F;
			14'd8340: ff_rdata <= 8'hFB;
			14'd8341: ff_rdata <= 8'hE6;
			14'd8342: ff_rdata <= 8'h7F;
			14'd8343: ff_rdata <= 8'h2A;
			14'd8344: ff_rdata <= 8'h95;
			14'd8345: ff_rdata <= 8'hF9;
			14'd8346: ff_rdata <= 8'hB5;
			14'd8347: ff_rdata <= 8'hB4;
			14'd8348: ff_rdata <= 8'h21;
			14'd8349: ff_rdata <= 8'h97;
			14'd8350: ff_rdata <= 8'hF9;
			14'd8351: ff_rdata <= 8'hB6;
			14'd8352: ff_rdata <= 8'hC4;
			14'd8353: ff_rdata <= 8'h8D;
			14'd8354: ff_rdata <= 8'h65;
			14'd8355: ff_rdata <= 8'hC9;
			14'd8356: ff_rdata <= 8'hED;
			14'd8357: ff_rdata <= 8'h4B;
			14'd8358: ff_rdata <= 8'h95;
			14'd8359: ff_rdata <= 8'hF9;
			14'd8360: ff_rdata <= 8'h78;
			14'd8361: ff_rdata <= 8'hB1;
			14'd8362: ff_rdata <= 8'h28;
			14'd8363: ff_rdata <= 8'h1E;
			14'd8364: ff_rdata <= 8'h69;
			14'd8365: ff_rdata <= 8'h60;
			14'd8366: ff_rdata <= 8'h3A;
			14'd8367: ff_rdata <= 8'h91;
			14'd8368: ff_rdata <= 8'hF9;
			14'd8369: ff_rdata <= 8'h47;
			14'd8370: ff_rdata <= 8'h3E;
			14'd8371: ff_rdata <= 8'h10;
			14'd8372: ff_rdata <= 8'h90;
			14'd8373: ff_rdata <= 8'h47;
			14'd8374: ff_rdata <= 8'h29;
			14'd8375: ff_rdata <= 8'h10;
			14'd8376: ff_rdata <= 8'hFD;
			14'd8377: ff_rdata <= 8'h3A;
			14'd8378: ff_rdata <= 8'h91;
			14'd8379: ff_rdata <= 8'hF9;
			14'd8380: ff_rdata <= 8'h3D;
			14'd8381: ff_rdata <= 8'hFA;
			14'd8382: ff_rdata <= 8'hCA;
			14'd8383: ff_rdata <= 8'h60;
			14'd8384: ff_rdata <= 8'h29;
			14'd8385: ff_rdata <= 8'hF5;
			14'd8386: ff_rdata <= 8'hE5;
			14'd8387: ff_rdata <= 8'hDC;
			14'd8388: ff_rdata <= 8'hCB;
			14'd8389: ff_rdata <= 8'h60;
			14'd8390: ff_rdata <= 8'hE1;
			14'd8391: ff_rdata <= 8'hF1;
			14'd8392: ff_rdata <= 8'h18;
			14'd8393: ff_rdata <= 8'hF2;
			14'd8394: ff_rdata <= 8'hC9;
			14'd8395: ff_rdata <= 8'h32;
			14'd8396: ff_rdata <= 8'h9A;
			14'd8397: ff_rdata <= 8'hF9;
			14'd8398: ff_rdata <= 8'hF3;
			14'd8399: ff_rdata <= 8'h2E;
			14'd8400: ff_rdata <= 8'h00;
			14'd8401: ff_rdata <= 8'hCD;
			14'd8402: ff_rdata <= 8'hE7;
			14'd8403: ff_rdata <= 8'h67;
			14'd8404: ff_rdata <= 8'h5E;
			14'd8405: ff_rdata <= 8'h23;
			14'd8406: ff_rdata <= 8'h56;
			14'd8407: ff_rdata <= 8'h7A;
			14'd8408: ff_rdata <= 8'hB3;
			14'd8409: ff_rdata <= 8'h28;
			14'd8410: ff_rdata <= 8'h08;
			14'd8411: ff_rdata <= 8'h1B;
			14'd8412: ff_rdata <= 8'h72;
			14'd8413: ff_rdata <= 8'h2B;
			14'd8414: ff_rdata <= 8'h73;
			14'd8415: ff_rdata <= 8'h7A;
			14'd8416: ff_rdata <= 8'hB3;
			14'd8417: ff_rdata <= 8'hC0;
			14'd8418: ff_rdata <= 8'h23;
			14'd8419: ff_rdata <= 8'h3A;
			14'd8420: ff_rdata <= 8'h92;
			14'd8421: ff_rdata <= 8'hF9;
			14'd8422: ff_rdata <= 8'h47;
			14'd8423: ff_rdata <= 8'h3A;
			14'd8424: ff_rdata <= 8'h9A;
			14'd8425: ff_rdata <= 8'hF9;
			14'd8426: ff_rdata <= 8'hB8;
			14'd8427: ff_rdata <= 8'hD2;
			14'd8428: ff_rdata <= 8'hFC;
			14'd8429: ff_rdata <= 8'h63;
			14'd8430: ff_rdata <= 8'hCD;
			14'd8431: ff_rdata <= 8'h88;
			14'd8432: ff_rdata <= 8'h63;
			14'd8433: ff_rdata <= 8'hC8;
			14'd8434: ff_rdata <= 8'h3C;
			14'd8435: ff_rdata <= 8'hCA;
			14'd8436: ff_rdata <= 8'h08;
			14'd8437: ff_rdata <= 8'h62;
			14'd8438: ff_rdata <= 8'h3D;
			14'd8439: ff_rdata <= 8'hFA;
			14'd8440: ff_rdata <= 8'h35;
			14'd8441: ff_rdata <= 8'h62;
			14'd8442: ff_rdata <= 8'hE5;
			14'd8443: ff_rdata <= 8'h57;
			14'd8444: ff_rdata <= 8'h5F;
			14'd8445: ff_rdata <= 8'h28;
			14'd8446: ff_rdata <= 8'h04;
			14'd8447: ff_rdata <= 8'hCD;
			14'd8448: ff_rdata <= 8'h88;
			14'd8449: ff_rdata <= 8'h63;
			14'd8450: ff_rdata <= 8'h5F;
			14'd8451: ff_rdata <= 8'h2E;
			14'd8452: ff_rdata <= 8'h0D;
			14'd8453: ff_rdata <= 8'hCD;
			14'd8454: ff_rdata <= 8'h96;
			14'd8455: ff_rdata <= 8'h63;
			14'd8456: ff_rdata <= 8'h73;
			14'd8457: ff_rdata <= 8'h23;
			14'd8458: ff_rdata <= 8'h72;
			14'd8459: ff_rdata <= 8'hE1;
			14'd8460: ff_rdata <= 8'hCD;
			14'd8461: ff_rdata <= 8'h88;
			14'd8462: ff_rdata <= 8'h63;
			14'd8463: ff_rdata <= 8'h4F;
			14'd8464: ff_rdata <= 8'hCD;
			14'd8465: ff_rdata <= 8'h88;
			14'd8466: ff_rdata <= 8'h63;
			14'd8467: ff_rdata <= 8'h77;
			14'd8468: ff_rdata <= 8'h2B;
			14'd8469: ff_rdata <= 8'h71;
			14'd8470: ff_rdata <= 8'h7A;
			14'd8471: ff_rdata <= 8'hB7;
			14'd8472: ff_rdata <= 8'hCA;
			14'd8473: ff_rdata <= 8'h77;
			14'd8474: ff_rdata <= 8'h61;
			14'd8475: ff_rdata <= 8'hCD;
			14'd8476: ff_rdata <= 8'hDA;
			14'd8477: ff_rdata <= 8'h61;
			14'd8478: ff_rdata <= 8'h2E;
			14'd8479: ff_rdata <= 8'h12;
			14'd8480: ff_rdata <= 8'hCD;
			14'd8481: ff_rdata <= 8'h96;
			14'd8482: ff_rdata <= 8'h63;
			14'd8483: ff_rdata <= 8'h4E;
			14'd8484: ff_rdata <= 8'hCD;
			14'd8485: ff_rdata <= 8'h3F;
			14'd8486: ff_rdata <= 8'h61;
			14'd8487: ff_rdata <= 8'hC2;
			14'd8488: ff_rdata <= 8'hBD;
			14'd8489: ff_rdata <= 8'h63;
			14'd8490: ff_rdata <= 8'hCD;
			14'd8491: ff_rdata <= 8'h9C;
			14'd8492: ff_rdata <= 8'h61;
			14'd8493: ff_rdata <= 8'hDA;
			14'd8494: ff_rdata <= 8'h72;
			14'd8495: ff_rdata <= 8'h61;
			14'd8496: ff_rdata <= 8'hC5;
			14'd8497: ff_rdata <= 8'hD5;
			14'd8498: ff_rdata <= 8'hCD;
			14'd8499: ff_rdata <= 8'h4A;
			14'd8500: ff_rdata <= 8'h6A;
			14'd8501: ff_rdata <= 8'h01;
			14'd8502: ff_rdata <= 8'h10;
			14'd8503: ff_rdata <= 8'h00;
			14'd8504: ff_rdata <= 8'hDD;
			14'd8505: ff_rdata <= 8'h09;
			14'd8506: ff_rdata <= 8'hD1;
			14'd8507: ff_rdata <= 8'hC1;
			14'd8508: ff_rdata <= 8'h10;
			14'd8509: ff_rdata <= 8'hF2;
			14'd8510: ff_rdata <= 8'hC9;
			14'd8511: ff_rdata <= 8'hE5;
			14'd8512: ff_rdata <= 8'h21;
			14'd8513: ff_rdata <= 8'h81;
			14'd8514: ff_rdata <= 8'hF9;
			14'd8515: ff_rdata <= 8'hCB;
			14'd8516: ff_rdata <= 8'h46;
			14'd8517: ff_rdata <= 8'hE1;
			14'd8518: ff_rdata <= 8'hC9;
			14'd8519: ff_rdata <= 8'hCD;
			14'd8520: ff_rdata <= 8'h88;
			14'd8521: ff_rdata <= 8'h63;
			14'd8522: ff_rdata <= 8'hC8;
			14'd8523: ff_rdata <= 8'hB7;
			14'd8524: ff_rdata <= 8'hFA;
			14'd8525: ff_rdata <= 8'hF2;
			14'd8526: ff_rdata <= 8'h60;
			14'd8527: ff_rdata <= 8'h28;
			14'd8528: ff_rdata <= 8'hA1;
			14'd8529: ff_rdata <= 8'h57;
			14'd8530: ff_rdata <= 8'hCD;
			14'd8531: ff_rdata <= 8'h88;
			14'd8532: ff_rdata <= 8'h63;
			14'd8533: ff_rdata <= 8'h5F;
			14'd8534: ff_rdata <= 8'hE5;
			14'd8535: ff_rdata <= 8'h2E;
			14'd8536: ff_rdata <= 8'h0D;
			14'd8537: ff_rdata <= 8'hCD;
			14'd8538: ff_rdata <= 8'h96;
			14'd8539: ff_rdata <= 8'h63;
			14'd8540: ff_rdata <= 8'h7B;
			14'd8541: ff_rdata <= 8'hBE;
			14'd8542: ff_rdata <= 8'h20;
			14'd8543: ff_rdata <= 8'h03;
			14'd8544: ff_rdata <= 8'h23;
			14'd8545: ff_rdata <= 8'h7A;
			14'd8546: ff_rdata <= 8'hBE;
			14'd8547: ff_rdata <= 8'hC2;
			14'd8548: ff_rdata <= 8'h03;
			14'd8549: ff_rdata <= 8'h61;
			14'd8550: ff_rdata <= 8'hE1;
			14'd8551: ff_rdata <= 8'hCD;
			14'd8552: ff_rdata <= 8'h88;
			14'd8553: ff_rdata <= 8'h63;
			14'd8554: ff_rdata <= 8'h4F;
			14'd8555: ff_rdata <= 8'hCD;
			14'd8556: ff_rdata <= 8'h88;
			14'd8557: ff_rdata <= 8'h63;
			14'd8558: ff_rdata <= 8'h77;
			14'd8559: ff_rdata <= 8'h2B;
			14'd8560: ff_rdata <= 8'h71;
			14'd8561: ff_rdata <= 8'hC9;
			14'd8562: ff_rdata <= 8'h3A;
			14'd8563: ff_rdata <= 8'h82;
			14'd8564: ff_rdata <= 8'hF9;
			14'd8565: ff_rdata <= 8'hC9;
			14'd8566: ff_rdata <= 8'hC9;
			14'd8567: ff_rdata <= 8'hCD;
			14'd8568: ff_rdata <= 8'h9C;
			14'd8569: ff_rdata <= 8'h61;
			14'd8570: ff_rdata <= 8'h30;
			14'd8571: ff_rdata <= 8'h0A;
			14'd8572: ff_rdata <= 8'hC0;
			14'd8573: ff_rdata <= 8'hCD;
			14'd8574: ff_rdata <= 8'h3F;
			14'd8575: ff_rdata <= 8'h61;
			14'd8576: ff_rdata <= 8'hC2;
			14'd8577: ff_rdata <= 8'hC8;
			14'd8578: ff_rdata <= 8'h63;
			14'd8579: ff_rdata <= 8'hC3;
			14'd8580: ff_rdata <= 8'h76;
			14'd8581: ff_rdata <= 8'h61;
			14'd8582: ff_rdata <= 8'hCD;
			14'd8583: ff_rdata <= 8'h3F;
			14'd8584: ff_rdata <= 8'h61;
			14'd8585: ff_rdata <= 8'hC2;
			14'd8586: ff_rdata <= 8'hC8;
			14'd8587: ff_rdata <= 8'h63;
			14'd8588: ff_rdata <= 8'hCD;
			14'd8589: ff_rdata <= 8'hDA;
			14'd8590: ff_rdata <= 8'h61;
			14'd8591: ff_rdata <= 8'hC5;
			14'd8592: ff_rdata <= 8'hCD;
			14'd8593: ff_rdata <= 8'h58;
			14'd8594: ff_rdata <= 8'h6C;
			14'd8595: ff_rdata <= 8'h01;
			14'd8596: ff_rdata <= 8'h10;
			14'd8597: ff_rdata <= 8'h00;
			14'd8598: ff_rdata <= 8'hDD;
			14'd8599: ff_rdata <= 8'h09;
			14'd8600: ff_rdata <= 8'hC1;
			14'd8601: ff_rdata <= 8'h10;
			14'd8602: ff_rdata <= 8'hF4;
			14'd8603: ff_rdata <= 8'hC9;
			14'd8604: ff_rdata <= 8'h3A;
			14'd8605: ff_rdata <= 8'h9A;
			14'd8606: ff_rdata <= 8'hF9;
			14'd8607: ff_rdata <= 8'h21;
			14'd8608: ff_rdata <= 8'h84;
			14'd8609: ff_rdata <= 8'hF9;
			14'd8610: ff_rdata <= 8'hBE;
			14'd8611: ff_rdata <= 8'h3F;
			14'd8612: ff_rdata <= 8'hD0;
			14'd8613: ff_rdata <= 8'hF5;
			14'd8614: ff_rdata <= 8'h3A;
			14'd8615: ff_rdata <= 8'h8E;
			14'd8616: ff_rdata <= 8'hF9;
			14'd8617: ff_rdata <= 8'h3D;
			14'd8618: ff_rdata <= 8'h28;
			14'd8619: ff_rdata <= 8'h02;
			14'd8620: ff_rdata <= 8'hF1;
			14'd8621: ff_rdata <= 8'hC9;
			14'd8622: ff_rdata <= 8'hF1;
			14'd8623: ff_rdata <= 8'h8F;
			14'd8624: ff_rdata <= 8'h1F;
			14'd8625: ff_rdata <= 8'hC9;
			14'd8626: ff_rdata <= 8'hCD;
			14'd8627: ff_rdata <= 8'h3F;
			14'd8628: ff_rdata <= 8'h61;
			14'd8629: ff_rdata <= 8'hC2;
			14'd8630: ff_rdata <= 8'hCC;
			14'd8631: ff_rdata <= 8'h63;
			14'd8632: ff_rdata <= 8'hCD;
			14'd8633: ff_rdata <= 8'h9C;
			14'd8634: ff_rdata <= 8'h61;
			14'd8635: ff_rdata <= 8'h30;
			14'd8636: ff_rdata <= 8'h05;
			14'd8637: ff_rdata <= 8'h79;
			14'd8638: ff_rdata <= 8'h32;
			14'd8639: ff_rdata <= 8'h82;
			14'd8640: ff_rdata <= 8'hF9;
			14'd8641: ff_rdata <= 8'hC9;
			14'd8642: ff_rdata <= 8'hC5;
			14'd8643: ff_rdata <= 8'hCD;
			14'd8644: ff_rdata <= 8'hDA;
			14'd8645: ff_rdata <= 8'h61;
			14'd8646: ff_rdata <= 8'hD1;
			14'd8647: ff_rdata <= 8'h4B;
			14'd8648: ff_rdata <= 8'hC5;
			14'd8649: ff_rdata <= 8'hCD;
			14'd8650: ff_rdata <= 8'h47;
			14'd8651: ff_rdata <= 8'h6A;
			14'd8652: ff_rdata <= 8'hC1;
			14'd8653: ff_rdata <= 8'hC5;
			14'd8654: ff_rdata <= 8'hCD;
			14'd8655: ff_rdata <= 8'hE1;
			14'd8656: ff_rdata <= 8'h68;
			14'd8657: ff_rdata <= 8'h01;
			14'd8658: ff_rdata <= 8'h10;
			14'd8659: ff_rdata <= 8'h00;
			14'd8660: ff_rdata <= 8'hDD;
			14'd8661: ff_rdata <= 8'h09;
			14'd8662: ff_rdata <= 8'hC1;
			14'd8663: ff_rdata <= 8'h10;
			14'd8664: ff_rdata <= 8'hEF;
			14'd8665: ff_rdata <= 8'hC9;
			14'd8666: ff_rdata <= 8'h3A;
			14'd8667: ff_rdata <= 8'h9A;
			14'd8668: ff_rdata <= 8'hF9;
			14'd8669: ff_rdata <= 8'hCD;
			14'd8670: ff_rdata <= 8'h9F;
			14'd8671: ff_rdata <= 8'h61;
			14'd8672: ff_rdata <= 8'h30;
			14'd8673: ff_rdata <= 8'h09;
			14'd8674: ff_rdata <= 8'h28;
			14'd8675: ff_rdata <= 8'h07;
			14'd8676: ff_rdata <= 8'hDD;
			14'd8677: ff_rdata <= 8'h21;
			14'd8678: ff_rdata <= 8'h87;
			14'd8679: ff_rdata <= 8'hFA;
			14'd8680: ff_rdata <= 8'h06;
			14'd8681: ff_rdata <= 8'h03;
			14'd8682: ff_rdata <= 8'hC9;
			14'd8683: ff_rdata <= 8'h21;
			14'd8684: ff_rdata <= 8'h85;
			14'd8685: ff_rdata <= 8'hF9;
			14'd8686: ff_rdata <= 8'hB7;
			14'd8687: ff_rdata <= 8'h28;
			14'd8688: ff_rdata <= 8'h06;
			14'd8689: ff_rdata <= 8'h47;
			14'd8690: ff_rdata <= 8'hAF;
			14'd8691: ff_rdata <= 8'h86;
			14'd8692: ff_rdata <= 8'h23;
			14'd8693: ff_rdata <= 8'h10;
			14'd8694: ff_rdata <= 8'hFC;
			14'd8695: ff_rdata <= 8'hDD;
			14'd8696: ff_rdata <= 8'h21;
			14'd8697: ff_rdata <= 8'h27;
			14'd8698: ff_rdata <= 8'hFA;
			14'd8699: ff_rdata <= 8'hB7;
			14'd8700: ff_rdata <= 8'h28;
			14'd8701: ff_rdata <= 8'h08;
			14'd8702: ff_rdata <= 8'h01;
			14'd8703: ff_rdata <= 8'h10;
			14'd8704: ff_rdata <= 8'h00;
			14'd8705: ff_rdata <= 8'hDD;
			14'd8706: ff_rdata <= 8'h09;
			14'd8707: ff_rdata <= 8'h3D;
			14'd8708: ff_rdata <= 8'h20;
			14'd8709: ff_rdata <= 8'hFB;
			14'd8710: ff_rdata <= 8'h46;
			14'd8711: ff_rdata <= 8'hC9;
			14'd8712: ff_rdata <= 8'hCD;
			14'd8713: ff_rdata <= 8'h77;
			14'd8714: ff_rdata <= 8'h61;
			14'd8715: ff_rdata <= 8'h2E;
			14'd8716: ff_rdata <= 8'h0D;
			14'd8717: ff_rdata <= 8'hCD;
			14'd8718: ff_rdata <= 8'h96;
			14'd8719: ff_rdata <= 8'h63;
			14'd8720: ff_rdata <= 8'h36;
			14'd8721: ff_rdata <= 8'h00;
			14'd8722: ff_rdata <= 8'h23;
			14'd8723: ff_rdata <= 8'h36;
			14'd8724: ff_rdata <= 8'h00;
			14'd8725: ff_rdata <= 8'h3A;
			14'd8726: ff_rdata <= 8'h9A;
			14'd8727: ff_rdata <= 8'hF9;
			14'd8728: ff_rdata <= 8'h21;
			14'd8729: ff_rdata <= 8'h01;
			14'd8730: ff_rdata <= 8'h00;
			14'd8731: ff_rdata <= 8'h47;
			14'd8732: ff_rdata <= 8'hB7;
			14'd8733: ff_rdata <= 8'h28;
			14'd8734: ff_rdata <= 8'h03;
			14'd8735: ff_rdata <= 8'h29;
			14'd8736: ff_rdata <= 8'h10;
			14'd8737: ff_rdata <= 8'hFD;
			14'd8738: ff_rdata <= 8'hEB;
			14'd8739: ff_rdata <= 8'hF3;
			14'd8740: ff_rdata <= 8'h2A;
			14'd8741: ff_rdata <= 8'h95;
			14'd8742: ff_rdata <= 8'hF9;
			14'd8743: ff_rdata <= 8'h7B;
			14'd8744: ff_rdata <= 8'hA5;
			14'd8745: ff_rdata <= 8'hAD;
			14'd8746: ff_rdata <= 8'h6F;
			14'd8747: ff_rdata <= 8'h7A;
			14'd8748: ff_rdata <= 8'hA4;
			14'd8749: ff_rdata <= 8'hAC;
			14'd8750: ff_rdata <= 8'h67;
			14'd8751: ff_rdata <= 8'h22;
			14'd8752: ff_rdata <= 8'h95;
			14'd8753: ff_rdata <= 8'hF9;
			14'd8754: ff_rdata <= 8'hC3;
			14'd8755: ff_rdata <= 8'h3D;
			14'd8756: ff_rdata <= 8'h68;
			14'd8757: ff_rdata <= 8'h5F;
			14'd8758: ff_rdata <= 8'hE6;
			14'd8759: ff_rdata <= 8'hC0;
			14'd8760: ff_rdata <= 8'hFE;
			14'd8761: ff_rdata <= 8'hC0;
			14'd8762: ff_rdata <= 8'hCA;
			14'd8763: ff_rdata <= 8'h41;
			14'd8764: ff_rdata <= 8'h63;
			14'd8765: ff_rdata <= 8'h7B;
			14'd8766: ff_rdata <= 8'h87;
			14'd8767: ff_rdata <= 8'hEB;
			14'd8768: ff_rdata <= 8'hC6;
			14'd8769: ff_rdata <= 8'h4E;
			14'd8770: ff_rdata <= 8'h6F;
			14'd8771: ff_rdata <= 8'h3E;
			14'd8772: ff_rdata <= 8'h00;
			14'd8773: ff_rdata <= 8'hCE;
			14'd8774: ff_rdata <= 8'h62;
			14'd8775: ff_rdata <= 8'h67;
			14'd8776: ff_rdata <= 8'h4E;
			14'd8777: ff_rdata <= 8'h23;
			14'd8778: ff_rdata <= 8'h46;
			14'd8779: ff_rdata <= 8'hEB;
			14'd8780: ff_rdata <= 8'hC5;
			14'd8781: ff_rdata <= 8'hC9;
			14'd8782: ff_rdata <= 8'h6E;
			14'd8783: ff_rdata <= 8'h62;
			14'd8784: ff_rdata <= 8'h71;
			14'd8785: ff_rdata <= 8'h62;
			14'd8786: ff_rdata <= 8'h9E;
			14'd8787: ff_rdata <= 8'h62;
			14'd8788: ff_rdata <= 8'hAC;
			14'd8789: ff_rdata <= 8'h62;
			14'd8790: ff_rdata <= 8'hB7;
			14'd8791: ff_rdata <= 8'h62;
			14'd8792: ff_rdata <= 8'hC1;
			14'd8793: ff_rdata <= 8'h62;
			14'd8794: ff_rdata <= 8'h18;
			14'd8795: ff_rdata <= 8'h63;
			14'd8796: ff_rdata <= 8'h47;
			14'd8797: ff_rdata <= 8'h61;
			14'd8798: ff_rdata <= 8'h64;
			14'd8799: ff_rdata <= 8'h62;
			14'd8800: ff_rdata <= 8'h66;
			14'd8801: ff_rdata <= 8'h62;
			14'd8802: ff_rdata <= 8'hF4;
			14'd8803: ff_rdata <= 8'h63;
			14'd8804: ff_rdata <= 8'hAF;
			14'd8805: ff_rdata <= 8'h01;
			14'd8806: ff_rdata <= 8'h3E;
			14'd8807: ff_rdata <= 8'h01;
			14'd8808: ff_rdata <= 8'h32;
			14'd8809: ff_rdata <= 8'h81;
			14'd8810: ff_rdata <= 8'hF9;
			14'd8811: ff_rdata <= 8'hC3;
			14'd8812: ff_rdata <= 8'hEE;
			14'd8813: ff_rdata <= 8'h60;
			14'd8814: ff_rdata <= 8'hC3;
			14'd8815: ff_rdata <= 8'h77;
			14'd8816: ff_rdata <= 8'h61;
			14'd8817: ff_rdata <= 8'hE5;
			14'd8818: ff_rdata <= 8'hCD;
			14'd8819: ff_rdata <= 8'h9C;
			14'd8820: ff_rdata <= 8'h61;
			14'd8821: ff_rdata <= 8'hE1;
			14'd8822: ff_rdata <= 8'h30;
			14'd8823: ff_rdata <= 8'h05;
			14'd8824: ff_rdata <= 8'hC2;
			14'd8825: ff_rdata <= 8'h00;
			14'd8826: ff_rdata <= 8'h63;
			14'd8827: ff_rdata <= 8'h18;
			14'd8828: ff_rdata <= 8'h0E;
			14'd8829: ff_rdata <= 8'hE5;
			14'd8830: ff_rdata <= 8'h2E;
			14'd8831: ff_rdata <= 8'h12;
			14'd8832: ff_rdata <= 8'hCD;
			14'd8833: ff_rdata <= 8'h96;
			14'd8834: ff_rdata <= 8'h63;
			14'd8835: ff_rdata <= 8'hCD;
			14'd8836: ff_rdata <= 8'h88;
			14'd8837: ff_rdata <= 8'h63;
			14'd8838: ff_rdata <= 8'h77;
			14'd8839: ff_rdata <= 8'hE1;
			14'd8840: ff_rdata <= 8'hC3;
			14'd8841: ff_rdata <= 8'hEE;
			14'd8842: ff_rdata <= 8'h60;
			14'd8843: ff_rdata <= 8'hE5;
			14'd8844: ff_rdata <= 8'h2E;
			14'd8845: ff_rdata <= 8'h12;
			14'd8846: ff_rdata <= 8'hCD;
			14'd8847: ff_rdata <= 8'h96;
			14'd8848: ff_rdata <= 8'h63;
			14'd8849: ff_rdata <= 8'hCD;
			14'd8850: ff_rdata <= 8'h88;
			14'd8851: ff_rdata <= 8'h63;
			14'd8852: ff_rdata <= 8'h77;
			14'd8853: ff_rdata <= 8'h87;
			14'd8854: ff_rdata <= 8'h87;
			14'd8855: ff_rdata <= 8'hC6;
			14'd8856: ff_rdata <= 8'h03;
			14'd8857: ff_rdata <= 8'hCD;
			14'd8858: ff_rdata <= 8'hF9;
			14'd8859: ff_rdata <= 8'h62;
			14'd8860: ff_rdata <= 8'h18;
			14'd8861: ff_rdata <= 8'hE9;
			14'd8862: ff_rdata <= 8'hE5;
			14'd8863: ff_rdata <= 8'hCD;
			14'd8864: ff_rdata <= 8'h88;
			14'd8865: ff_rdata <= 8'h63;
			14'd8866: ff_rdata <= 8'h4F;
			14'd8867: ff_rdata <= 8'hCD;
			14'd8868: ff_rdata <= 8'h88;
			14'd8869: ff_rdata <= 8'h63;
			14'd8870: ff_rdata <= 8'h47;
			14'd8871: ff_rdata <= 8'hCD;
			14'd8872: ff_rdata <= 8'hB5;
			14'd8873: ff_rdata <= 8'h6D;
			14'd8874: ff_rdata <= 8'h18;
			14'd8875: ff_rdata <= 8'hDB;
			14'd8876: ff_rdata <= 8'hCD;
			14'd8877: ff_rdata <= 8'h88;
			14'd8878: ff_rdata <= 8'h63;
			14'd8879: ff_rdata <= 8'h4F;
			14'd8880: ff_rdata <= 8'hCD;
			14'd8881: ff_rdata <= 8'h88;
			14'd8882: ff_rdata <= 8'h63;
			14'd8883: ff_rdata <= 8'h77;
			14'd8884: ff_rdata <= 8'h2B;
			14'd8885: ff_rdata <= 8'h71;
			14'd8886: ff_rdata <= 8'hC9;
			14'd8887: ff_rdata <= 8'hE5;
			14'd8888: ff_rdata <= 8'hCD;
			14'd8889: ff_rdata <= 8'h88;
			14'd8890: ff_rdata <= 8'h63;
			14'd8891: ff_rdata <= 8'h4F;
			14'd8892: ff_rdata <= 8'hCD;
			14'd8893: ff_rdata <= 8'hB2;
			14'd8894: ff_rdata <= 8'h61;
			14'd8895: ff_rdata <= 8'h18;
			14'd8896: ff_rdata <= 8'hC6;
			14'd8897: ff_rdata <= 8'hCD;
			14'd8898: ff_rdata <= 8'h3F;
			14'd8899: ff_rdata <= 8'h61;
			14'd8900: ff_rdata <= 8'hC2;
			14'd8901: ff_rdata <= 8'hD1;
			14'd8902: ff_rdata <= 8'h63;
			14'd8903: ff_rdata <= 8'hE5;
			14'd8904: ff_rdata <= 8'hCD;
			14'd8905: ff_rdata <= 8'h9C;
			14'd8906: ff_rdata <= 8'h61;
			14'd8907: ff_rdata <= 8'h30;
			14'd8908: ff_rdata <= 8'h09;
			14'd8909: ff_rdata <= 8'h28;
			14'd8910: ff_rdata <= 8'h1E;
			14'd8911: ff_rdata <= 8'hCD;
			14'd8912: ff_rdata <= 8'hDA;
			14'd8913: ff_rdata <= 8'h61;
			14'd8914: ff_rdata <= 8'h06;
			14'd8915: ff_rdata <= 8'h01;
			14'd8916: ff_rdata <= 8'h18;
			14'd8917: ff_rdata <= 8'h03;
			14'd8918: ff_rdata <= 8'hCD;
			14'd8919: ff_rdata <= 8'hDA;
			14'd8920: ff_rdata <= 8'h61;
			14'd8921: ff_rdata <= 8'hCD;
			14'd8922: ff_rdata <= 8'h88;
			14'd8923: ff_rdata <= 8'h63;
			14'd8924: ff_rdata <= 8'h5F;
			14'd8925: ff_rdata <= 8'hC5;
			14'd8926: ff_rdata <= 8'hD5;
			14'd8927: ff_rdata <= 8'hCD;
			14'd8928: ff_rdata <= 8'hCC;
			14'd8929: ff_rdata <= 8'h69;
			14'd8930: ff_rdata <= 8'h01;
			14'd8931: ff_rdata <= 8'h10;
			14'd8932: ff_rdata <= 8'h00;
			14'd8933: ff_rdata <= 8'hDD;
			14'd8934: ff_rdata <= 8'h09;
			14'd8935: ff_rdata <= 8'hD1;
			14'd8936: ff_rdata <= 8'hC1;
			14'd8937: ff_rdata <= 8'h10;
			14'd8938: ff_rdata <= 8'hF2;
			14'd8939: ff_rdata <= 8'h18;
			14'd8940: ff_rdata <= 8'h9A;
			14'd8941: ff_rdata <= 8'hCD;
			14'd8942: ff_rdata <= 8'h88;
			14'd8943: ff_rdata <= 8'h63;
			14'd8944: ff_rdata <= 8'h5F;
			14'd8945: ff_rdata <= 8'h3E;
			14'd8946: ff_rdata <= 8'h3F;
			14'd8947: ff_rdata <= 8'h93;
			14'd8948: ff_rdata <= 8'hCD;
			14'd8949: ff_rdata <= 8'hF9;
			14'd8950: ff_rdata <= 8'h62;
			14'd8951: ff_rdata <= 8'hE1;
			14'd8952: ff_rdata <= 8'hC9;
			14'd8953: ff_rdata <= 8'h4F;
			14'd8954: ff_rdata <= 8'h06;
			14'd8955: ff_rdata <= 8'h00;
			14'd8956: ff_rdata <= 8'h5F;
			14'd8957: ff_rdata <= 8'h16;
			14'd8958: ff_rdata <= 8'h00;
			14'd8959: ff_rdata <= 8'hC9;
			14'd8960: ff_rdata <= 8'hE5;
			14'd8961: ff_rdata <= 8'h2E;
			14'd8962: ff_rdata <= 8'h0A;
			14'd8963: ff_rdata <= 8'hCD;
			14'd8964: ff_rdata <= 8'h96;
			14'd8965: ff_rdata <= 8'h63;
			14'd8966: ff_rdata <= 8'hCD;
			14'd8967: ff_rdata <= 8'h88;
			14'd8968: ff_rdata <= 8'h63;
			14'd8969: ff_rdata <= 8'h77;
			14'd8970: ff_rdata <= 8'h5F;
			14'd8971: ff_rdata <= 8'h2E;
			14'd8972: ff_rdata <= 8'h08;
			14'd8973: ff_rdata <= 8'hCD;
			14'd8974: ff_rdata <= 8'h96;
			14'd8975: ff_rdata <= 8'h63;
			14'd8976: ff_rdata <= 8'h7E;
			14'd8977: ff_rdata <= 8'h2F;
			14'd8978: ff_rdata <= 8'hCD;
			14'd8979: ff_rdata <= 8'h2F;
			14'd8980: ff_rdata <= 8'h63;
			14'd8981: ff_rdata <= 8'hC3;
			14'd8982: ff_rdata <= 8'h87;
			14'd8983: ff_rdata <= 8'h62;
			14'd8984: ff_rdata <= 8'hE5;
			14'd8985: ff_rdata <= 8'h2E;
			14'd8986: ff_rdata <= 8'h0C;
			14'd8987: ff_rdata <= 8'hCD;
			14'd8988: ff_rdata <= 8'h96;
			14'd8989: ff_rdata <= 8'h63;
			14'd8990: ff_rdata <= 8'hCD;
			14'd8991: ff_rdata <= 8'h88;
			14'd8992: ff_rdata <= 8'h63;
			14'd8993: ff_rdata <= 8'h77;
			14'd8994: ff_rdata <= 8'h5F;
			14'd8995: ff_rdata <= 8'h2E;
			14'd8996: ff_rdata <= 8'h08;
			14'd8997: ff_rdata <= 8'hCD;
			14'd8998: ff_rdata <= 8'h96;
			14'd8999: ff_rdata <= 8'h63;
			14'd9000: ff_rdata <= 8'h7E;
			14'd9001: ff_rdata <= 8'hCD;
			14'd9002: ff_rdata <= 8'h2F;
			14'd9003: ff_rdata <= 8'h63;
			14'd9004: ff_rdata <= 8'hC3;
			14'd9005: ff_rdata <= 8'h87;
			14'd9006: ff_rdata <= 8'h62;
			14'd9007: ff_rdata <= 8'hE6;
			14'd9008: ff_rdata <= 8'h1F;
			14'd9009: ff_rdata <= 8'hC8;
			14'd9010: ff_rdata <= 8'hCD;
			14'd9011: ff_rdata <= 8'h3F;
			14'd9012: ff_rdata <= 8'h61;
			14'd9013: ff_rdata <= 8'hC2;
			14'd9014: ff_rdata <= 8'hE4;
			14'd9015: ff_rdata <= 8'h63;
			14'd9016: ff_rdata <= 8'hC5;
			14'd9017: ff_rdata <= 8'hD5;
			14'd9018: ff_rdata <= 8'h4F;
			14'd9019: ff_rdata <= 8'hCD;
			14'd9020: ff_rdata <= 8'hDB;
			14'd9021: ff_rdata <= 8'h69;
			14'd9022: ff_rdata <= 8'hD1;
			14'd9023: ff_rdata <= 8'hC1;
			14'd9024: ff_rdata <= 8'hC9;
			14'd9025: ff_rdata <= 8'hCD;
			14'd9026: ff_rdata <= 8'h88;
			14'd9027: ff_rdata <= 8'h63;
			14'd9028: ff_rdata <= 8'h57;
			14'd9029: ff_rdata <= 8'hCD;
			14'd9030: ff_rdata <= 8'h88;
			14'd9031: ff_rdata <= 8'h63;
			14'd9032: ff_rdata <= 8'h4F;
			14'd9033: ff_rdata <= 8'hCD;
			14'd9034: ff_rdata <= 8'h88;
			14'd9035: ff_rdata <= 8'h63;
			14'd9036: ff_rdata <= 8'h77;
			14'd9037: ff_rdata <= 8'h2B;
			14'd9038: ff_rdata <= 8'h71;
			14'd9039: ff_rdata <= 8'hE5;
			14'd9040: ff_rdata <= 8'h2E;
			14'd9041: ff_rdata <= 8'h08;
			14'd9042: ff_rdata <= 8'hCD;
			14'd9043: ff_rdata <= 8'h96;
			14'd9044: ff_rdata <= 8'h63;
			14'd9045: ff_rdata <= 8'h7A;
			14'd9046: ff_rdata <= 8'hAE;
			14'd9047: ff_rdata <= 8'h28;
			14'd9048: ff_rdata <= 8'h20;
			14'd9049: ff_rdata <= 8'h72;
			14'd9050: ff_rdata <= 8'hD5;
			14'd9051: ff_rdata <= 8'hF5;
			14'd9052: ff_rdata <= 8'hA2;
			14'd9053: ff_rdata <= 8'hF5;
			14'd9054: ff_rdata <= 8'h2E;
			14'd9055: ff_rdata <= 8'h0C;
			14'd9056: ff_rdata <= 8'hCD;
			14'd9057: ff_rdata <= 8'h96;
			14'd9058: ff_rdata <= 8'h63;
			14'd9059: ff_rdata <= 8'h5E;
			14'd9060: ff_rdata <= 8'hF1;
			14'd9061: ff_rdata <= 8'hCD;
			14'd9062: ff_rdata <= 8'h2F;
			14'd9063: ff_rdata <= 8'h63;
			14'd9064: ff_rdata <= 8'h7A;
			14'd9065: ff_rdata <= 8'h2F;
			14'd9066: ff_rdata <= 8'h57;
			14'd9067: ff_rdata <= 8'hF1;
			14'd9068: ff_rdata <= 8'hA2;
			14'd9069: ff_rdata <= 8'hF5;
			14'd9070: ff_rdata <= 8'h2E;
			14'd9071: ff_rdata <= 8'h0A;
			14'd9072: ff_rdata <= 8'hCD;
			14'd9073: ff_rdata <= 8'h96;
			14'd9074: ff_rdata <= 8'h63;
			14'd9075: ff_rdata <= 8'h5E;
			14'd9076: ff_rdata <= 8'hF1;
			14'd9077: ff_rdata <= 8'hCD;
			14'd9078: ff_rdata <= 8'h2F;
			14'd9079: ff_rdata <= 8'h63;
			14'd9080: ff_rdata <= 8'hD1;
			14'd9081: ff_rdata <= 8'hE1;
			14'd9082: ff_rdata <= 8'h7B;
			14'd9083: ff_rdata <= 8'hE6;
			14'd9084: ff_rdata <= 8'h3F;
			14'd9085: ff_rdata <= 8'h4F;
			14'd9086: ff_rdata <= 8'hCD;
			14'd9087: ff_rdata <= 8'h3F;
			14'd9088: ff_rdata <= 8'h61;
			14'd9089: ff_rdata <= 8'hC2;
			14'd9090: ff_rdata <= 8'hEF;
			14'd9091: ff_rdata <= 8'h63;
			14'd9092: ff_rdata <= 8'hCD;
			14'd9093: ff_rdata <= 8'h68;
			14'd9094: ff_rdata <= 8'h6C;
			14'd9095: ff_rdata <= 8'hC9;
			14'd9096: ff_rdata <= 8'hE5;
			14'd9097: ff_rdata <= 8'hD5;
			14'd9098: ff_rdata <= 8'hC5;
			14'd9099: ff_rdata <= 8'h3A;
			14'd9100: ff_rdata <= 8'h9A;
			14'd9101: ff_rdata <= 8'hF9;
			14'd9102: ff_rdata <= 8'hF3;
			14'd9103: ff_rdata <= 8'hCD;
			14'd9104: ff_rdata <= 8'h14;
			14'd9105: ff_rdata <= 8'h67;
			14'd9106: ff_rdata <= 8'hC1;
			14'd9107: ff_rdata <= 8'hD1;
			14'd9108: ff_rdata <= 8'hE1;
			14'd9109: ff_rdata <= 8'hC9;
			14'd9110: ff_rdata <= 8'h3A;
			14'd9111: ff_rdata <= 8'h9A;
			14'd9112: ff_rdata <= 8'hF9;
			14'd9113: ff_rdata <= 8'hF3;
			14'd9114: ff_rdata <= 8'hC3;
			14'd9115: ff_rdata <= 8'hE7;
			14'd9116: ff_rdata <= 8'h67;
			14'd9117: ff_rdata <= 8'hFB;
			14'd9118: ff_rdata <= 8'hCD;
			14'd9119: ff_rdata <= 8'hB1;
			14'd9120: ff_rdata <= 8'h63;
			14'd9121: ff_rdata <= 8'h37;
			14'd9122: ff_rdata <= 8'hC8;
			14'd9123: ff_rdata <= 8'hF3;
			14'd9124: ff_rdata <= 8'h2A;
			14'd9125: ff_rdata <= 8'h95;
			14'd9126: ff_rdata <= 8'hF9;
			14'd9127: ff_rdata <= 8'h7D;
			14'd9128: ff_rdata <= 8'hB4;
			14'd9129: ff_rdata <= 8'h21;
			14'd9130: ff_rdata <= 8'h97;
			14'd9131: ff_rdata <= 8'hF9;
			14'd9132: ff_rdata <= 8'hB6;
			14'd9133: ff_rdata <= 8'h20;
			14'd9134: ff_rdata <= 8'hEE;
			14'd9135: ff_rdata <= 8'hFB;
			14'd9136: ff_rdata <= 8'hC9;
			14'd9137: ff_rdata <= 8'h3A;
			14'd9138: ff_rdata <= 8'hB1;
			14'd9139: ff_rdata <= 8'hFB;
			14'd9140: ff_rdata <= 8'hB7;
			14'd9141: ff_rdata <= 8'hC0;
			14'd9142: ff_rdata <= 8'h3A;
			14'd9143: ff_rdata <= 8'h9B;
			14'd9144: ff_rdata <= 8'hFC;
			14'd9145: ff_rdata <= 8'hD6;
			14'd9146: ff_rdata <= 8'h03;
			14'd9147: ff_rdata <= 8'hB7;
			14'd9148: ff_rdata <= 8'hC9;
			14'd9149: ff_rdata <= 8'h06;
			14'd9150: ff_rdata <= 8'h00;
			14'd9151: ff_rdata <= 8'h3A;
			14'd9152: ff_rdata <= 8'h9A;
			14'd9153: ff_rdata <= 8'hF9;
			14'd9154: ff_rdata <= 8'hE5;
			14'd9155: ff_rdata <= 8'hCD;
			14'd9156: ff_rdata <= 8'h75;
			14'd9157: ff_rdata <= 8'hF9;
			14'd9158: ff_rdata <= 8'hE1;
			14'd9159: ff_rdata <= 8'hC9;
			14'd9160: ff_rdata <= 8'h06;
			14'd9161: ff_rdata <= 8'h01;
			14'd9162: ff_rdata <= 8'h18;
			14'd9163: ff_rdata <= 8'hF3;
			14'd9164: ff_rdata <= 8'h06;
			14'd9165: ff_rdata <= 8'h02;
			14'd9166: ff_rdata <= 8'h51;
			14'd9167: ff_rdata <= 8'h18;
			14'd9168: ff_rdata <= 8'hEE;
			14'd9169: ff_rdata <= 8'hCD;
			14'd9170: ff_rdata <= 8'h88;
			14'd9171: ff_rdata <= 8'h63;
			14'd9172: ff_rdata <= 8'h57;
			14'd9173: ff_rdata <= 8'hE5;
			14'd9174: ff_rdata <= 8'hCD;
			14'd9175: ff_rdata <= 8'h9C;
			14'd9176: ff_rdata <= 8'h61;
			14'd9177: ff_rdata <= 8'hE1;
			14'd9178: ff_rdata <= 8'h06;
			14'd9179: ff_rdata <= 8'h03;
			14'd9180: ff_rdata <= 8'h30;
			14'd9181: ff_rdata <= 8'hE1;
			14'd9182: ff_rdata <= 8'h28;
			14'd9183: ff_rdata <= 8'hDF;
			14'd9184: ff_rdata <= 8'h06;
			14'd9185: ff_rdata <= 8'h04;
			14'd9186: ff_rdata <= 8'h18;
			14'd9187: ff_rdata <= 8'hDB;
			14'd9188: ff_rdata <= 8'hC5;
			14'd9189: ff_rdata <= 8'hD5;
			14'd9190: ff_rdata <= 8'h57;
			14'd9191: ff_rdata <= 8'h06;
			14'd9192: ff_rdata <= 8'h05;
			14'd9193: ff_rdata <= 8'hCD;
			14'd9194: ff_rdata <= 8'hBF;
			14'd9195: ff_rdata <= 8'h63;
			14'd9196: ff_rdata <= 8'hD1;
			14'd9197: ff_rdata <= 8'hC1;
			14'd9198: ff_rdata <= 8'hC9;
			14'd9199: ff_rdata <= 8'h06;
			14'd9200: ff_rdata <= 8'h06;
			14'd9201: ff_rdata <= 8'h51;
			14'd9202: ff_rdata <= 8'h18;
			14'd9203: ff_rdata <= 8'hCB;
			14'd9204: ff_rdata <= 8'hCD;
			14'd9205: ff_rdata <= 8'h88;
			14'd9206: ff_rdata <= 8'h63;
			14'd9207: ff_rdata <= 8'h57;
			14'd9208: ff_rdata <= 8'h06;
			14'd9209: ff_rdata <= 8'h07;
			14'd9210: ff_rdata <= 8'h18;
			14'd9211: ff_rdata <= 8'hC3;
			14'd9212: ff_rdata <= 8'h3A;
			14'd9213: ff_rdata <= 8'h92;
			14'd9214: ff_rdata <= 8'hF9;
			14'd9215: ff_rdata <= 8'h47;
			14'd9216: ff_rdata <= 8'h3A;
			14'd9217: ff_rdata <= 8'h9A;
			14'd9218: ff_rdata <= 8'hF9;
			14'd9219: ff_rdata <= 8'h90;
			14'd9220: ff_rdata <= 8'h47;
			14'd9221: ff_rdata <= 8'hCD;
			14'd9222: ff_rdata <= 8'h88;
			14'd9223: ff_rdata <= 8'h63;
			14'd9224: ff_rdata <= 8'hC8;
			14'd9225: ff_rdata <= 8'hFE;
			14'd9226: ff_rdata <= 8'hFF;
			14'd9227: ff_rdata <= 8'h28;
			14'd9228: ff_rdata <= 8'h5B;
			14'd9229: ff_rdata <= 8'h57;
			14'd9230: ff_rdata <= 8'hE6;
			14'd9231: ff_rdata <= 8'hE0;
			14'd9232: ff_rdata <= 8'h07;
			14'd9233: ff_rdata <= 8'h07;
			14'd9234: ff_rdata <= 8'h07;
			14'd9235: ff_rdata <= 8'h4F;
			14'd9236: ff_rdata <= 8'h7A;
			14'd9237: ff_rdata <= 8'hE6;
			14'd9238: ff_rdata <= 8'h1F;
			14'd9239: ff_rdata <= 8'h77;
			14'd9240: ff_rdata <= 8'hCD;
			14'd9241: ff_rdata <= 8'h88;
			14'd9242: ff_rdata <= 8'h63;
			14'd9243: ff_rdata <= 8'h2B;
			14'd9244: ff_rdata <= 8'h77;
			14'd9245: ff_rdata <= 8'h0C;
			14'd9246: ff_rdata <= 8'h0D;
			14'd9247: ff_rdata <= 8'hC8;
			14'd9248: ff_rdata <= 8'hCD;
			14'd9249: ff_rdata <= 8'h88;
			14'd9250: ff_rdata <= 8'h63;
			14'd9251: ff_rdata <= 8'h57;
			14'd9252: ff_rdata <= 8'hE6;
			14'd9253: ff_rdata <= 8'hC0;
			14'd9254: ff_rdata <= 8'h20;
			14'd9255: ff_rdata <= 8'h11;
			14'd9256: ff_rdata <= 8'hCD;
			14'd9257: ff_rdata <= 8'h88;
			14'd9258: ff_rdata <= 8'h63;
			14'd9259: ff_rdata <= 8'h5F;
			14'd9260: ff_rdata <= 8'h78;
			14'd9261: ff_rdata <= 8'h07;
			14'd9262: ff_rdata <= 8'hCD;
			14'd9263: ff_rdata <= 8'h80;
			14'd9264: ff_rdata <= 8'h64;
			14'd9265: ff_rdata <= 8'h3C;
			14'd9266: ff_rdata <= 8'h5A;
			14'd9267: ff_rdata <= 8'hCD;
			14'd9268: ff_rdata <= 8'h80;
			14'd9269: ff_rdata <= 8'h64;
			14'd9270: ff_rdata <= 8'h0D;
			14'd9271: ff_rdata <= 8'h18;
			14'd9272: ff_rdata <= 8'hE5;
			14'd9273: ff_rdata <= 8'h67;
			14'd9274: ff_rdata <= 8'hE6;
			14'd9275: ff_rdata <= 8'h80;
			14'd9276: ff_rdata <= 8'h28;
			14'd9277: ff_rdata <= 8'h0F;
			14'd9278: ff_rdata <= 8'h5A;
			14'd9279: ff_rdata <= 8'h78;
			14'd9280: ff_rdata <= 8'hC6;
			14'd9281: ff_rdata <= 8'h08;
			14'd9282: ff_rdata <= 8'hCD;
			14'd9283: ff_rdata <= 8'h80;
			14'd9284: ff_rdata <= 8'h64;
			14'd9285: ff_rdata <= 8'h7B;
			14'd9286: ff_rdata <= 8'hE6;
			14'd9287: ff_rdata <= 8'h10;
			14'd9288: ff_rdata <= 8'h3E;
			14'd9289: ff_rdata <= 8'h0D;
			14'd9290: ff_rdata <= 8'hC4;
			14'd9291: ff_rdata <= 8'h80;
			14'd9292: ff_rdata <= 8'h64;
			14'd9293: ff_rdata <= 8'h7C;
			14'd9294: ff_rdata <= 8'hE6;
			14'd9295: ff_rdata <= 8'h40;
			14'd9296: ff_rdata <= 8'h28;
			14'd9297: ff_rdata <= 8'hCC;
			14'd9298: ff_rdata <= 8'hCD;
			14'd9299: ff_rdata <= 8'h88;
			14'd9300: ff_rdata <= 8'h63;
			14'd9301: ff_rdata <= 8'h57;
			14'd9302: ff_rdata <= 8'hCD;
			14'd9303: ff_rdata <= 8'h88;
			14'd9304: ff_rdata <= 8'h63;
			14'd9305: ff_rdata <= 8'h5F;
			14'd9306: ff_rdata <= 8'h3E;
			14'd9307: ff_rdata <= 8'h0B;
			14'd9308: ff_rdata <= 8'hCD;
			14'd9309: ff_rdata <= 8'h80;
			14'd9310: ff_rdata <= 8'h64;
			14'd9311: ff_rdata <= 8'h3C;
			14'd9312: ff_rdata <= 8'h5A;
			14'd9313: ff_rdata <= 8'hCD;
			14'd9314: ff_rdata <= 8'h80;
			14'd9315: ff_rdata <= 8'h64;
			14'd9316: ff_rdata <= 8'h0D;
			14'd9317: ff_rdata <= 8'h0D;
			14'd9318: ff_rdata <= 8'h18;
			14'd9319: ff_rdata <= 8'hB6;
			14'd9320: ff_rdata <= 8'h78;
			14'd9321: ff_rdata <= 8'hC6;
			14'd9322: ff_rdata <= 8'h08;
			14'd9323: ff_rdata <= 8'h1E;
			14'd9324: ff_rdata <= 8'h00;
			14'd9325: ff_rdata <= 8'hCD;
			14'd9326: ff_rdata <= 8'h80;
			14'd9327: ff_rdata <= 8'h64;
			14'd9328: ff_rdata <= 8'h04;
			14'd9329: ff_rdata <= 8'hF3;
			14'd9330: ff_rdata <= 8'h21;
			14'd9331: ff_rdata <= 8'h3F;
			14'd9332: ff_rdata <= 8'hFB;
			14'd9333: ff_rdata <= 8'hAF;
			14'd9334: ff_rdata <= 8'h37;
			14'd9335: ff_rdata <= 8'h17;
			14'd9336: ff_rdata <= 8'h10;
			14'd9337: ff_rdata <= 8'hFD;
			14'd9338: ff_rdata <= 8'hA6;
			14'd9339: ff_rdata <= 8'hAE;
			14'd9340: ff_rdata <= 8'h77;
			14'd9341: ff_rdata <= 8'hC3;
			14'd9342: ff_rdata <= 8'h15;
			14'd9343: ff_rdata <= 8'h62;
			14'd9344: ff_rdata <= 8'hF3;
			14'd9345: ff_rdata <= 8'hD3;
			14'd9346: ff_rdata <= 8'hA0;
			14'd9347: ff_rdata <= 8'hF5;
			14'd9348: ff_rdata <= 8'h7B;
			14'd9349: ff_rdata <= 8'hD3;
			14'd9350: ff_rdata <= 8'hA1;
			14'd9351: ff_rdata <= 8'hF1;
			14'd9352: ff_rdata <= 8'hC9;
			14'd9353: ff_rdata <= 8'hAF;
			14'd9354: ff_rdata <= 8'h32;
			14'd9355: ff_rdata <= 8'h98;
			14'd9356: ff_rdata <= 8'hF9;
			14'd9357: ff_rdata <= 8'h3A;
			14'd9358: ff_rdata <= 8'h84;
			14'd9359: ff_rdata <= 8'hF9;
			14'd9360: ff_rdata <= 8'h21;
			14'd9361: ff_rdata <= 8'h8E;
			14'd9362: ff_rdata <= 8'hF9;
			14'd9363: ff_rdata <= 8'hCB;
			14'd9364: ff_rdata <= 8'h46;
			14'd9365: ff_rdata <= 8'h28;
			14'd9366: ff_rdata <= 8'h01;
			14'd9367: ff_rdata <= 8'h3C;
			14'd9368: ff_rdata <= 8'hCB;
			14'd9369: ff_rdata <= 8'h4E;
			14'd9370: ff_rdata <= 8'h28;
			14'd9371: ff_rdata <= 8'h01;
			14'd9372: ff_rdata <= 8'h3C;
			14'd9373: ff_rdata <= 8'h32;
			14'd9374: ff_rdata <= 8'h92;
			14'd9375: ff_rdata <= 8'hF9;
			14'd9376: ff_rdata <= 8'hC6;
			14'd9377: ff_rdata <= 8'h03;
			14'd9378: ff_rdata <= 8'h32;
			14'd9379: ff_rdata <= 8'h91;
			14'd9380: ff_rdata <= 8'hF9;
			14'd9381: ff_rdata <= 8'h47;
			14'd9382: ff_rdata <= 8'hF6;
			14'd9383: ff_rdata <= 8'h80;
			14'd9384: ff_rdata <= 8'h32;
			14'd9385: ff_rdata <= 8'h93;
			14'd9386: ff_rdata <= 8'hF9;
			14'd9387: ff_rdata <= 8'h21;
			14'd9388: ff_rdata <= 8'h00;
			14'd9389: ff_rdata <= 8'h00;
			14'd9390: ff_rdata <= 8'h37;
			14'd9391: ff_rdata <= 8'hED;
			14'd9392: ff_rdata <= 8'h6A;
			14'd9393: ff_rdata <= 8'h10;
			14'd9394: ff_rdata <= 8'hFB;
			14'd9395: ff_rdata <= 8'h22;
			14'd9396: ff_rdata <= 8'h8F;
			14'd9397: ff_rdata <= 8'hF9;
			14'd9398: ff_rdata <= 8'h3A;
			14'd9399: ff_rdata <= 8'h92;
			14'd9400: ff_rdata <= 8'hF9;
			14'd9401: ff_rdata <= 8'h21;
			14'd9402: ff_rdata <= 8'hE4;
			14'd9403: ff_rdata <= 8'h64;
			14'd9404: ff_rdata <= 8'hCD;
			14'd9405: ff_rdata <= 8'h86;
			14'd9406: ff_rdata <= 8'h54;
			14'd9407: ff_rdata <= 8'h7E;
			14'd9408: ff_rdata <= 8'h32;
			14'd9409: ff_rdata <= 8'h94;
			14'd9410: ff_rdata <= 8'hF9;
			14'd9411: ff_rdata <= 8'h2A;
			14'd9412: ff_rdata <= 8'h7D;
			14'd9413: ff_rdata <= 8'hF9;
			14'd9414: ff_rdata <= 8'h11;
			14'd9415: ff_rdata <= 8'h00;
			14'd9416: ff_rdata <= 8'h00;
			14'd9417: ff_rdata <= 8'h19;
			14'd9418: ff_rdata <= 8'h22;
			14'd9419: ff_rdata <= 8'h9B;
			14'd9420: ff_rdata <= 8'hF9;
			14'd9421: ff_rdata <= 8'h3A;
			14'd9422: ff_rdata <= 8'hC1;
			14'd9423: ff_rdata <= 8'hFC;
			14'd9424: ff_rdata <= 8'h21;
			14'd9425: ff_rdata <= 8'h2B;
			14'd9426: ff_rdata <= 8'h00;
			14'd9427: ff_rdata <= 8'hCD;
			14'd9428: ff_rdata <= 8'h0C;
			14'd9429: ff_rdata <= 8'h00;
			14'd9430: ff_rdata <= 8'hE6;
			14'd9431: ff_rdata <= 8'h80;
			14'd9432: ff_rdata <= 8'h21;
			14'd9433: ff_rdata <= 8'h40;
			14'd9434: ff_rdata <= 8'h38;
			14'd9435: ff_rdata <= 8'h28;
			14'd9436: ff_rdata <= 8'h03;
			14'd9437: ff_rdata <= 8'h21;
			14'd9438: ff_rdata <= 8'hE0;
			14'd9439: ff_rdata <= 8'h2E;
			14'd9440: ff_rdata <= 8'h22;
			14'd9441: ff_rdata <= 8'h7A;
			14'd9442: ff_rdata <= 8'hF9;
			14'd9443: ff_rdata <= 8'hC9;
			14'd9444: ff_rdata <= 8'h7F;
			14'd9445: ff_rdata <= 8'h3F;
			14'd9446: ff_rdata <= 8'h3F;
			14'd9447: ff_rdata <= 8'h3F;
			14'd9448: ff_rdata <= 8'h1F;
			14'd9449: ff_rdata <= 8'h1F;
			14'd9450: ff_rdata <= 8'h1F;
			14'd9451: ff_rdata <= 8'h1F;
			14'd9452: ff_rdata <= 8'h1F;
			14'd9453: ff_rdata <= 8'h1F;
			14'd9454: ff_rdata <= 8'hCD;
			14'd9455: ff_rdata <= 8'h89;
			14'd9456: ff_rdata <= 8'h67;
			14'd9457: ff_rdata <= 8'hF3;
			14'd9458: ff_rdata <= 8'hAF;
			14'd9459: ff_rdata <= 8'h32;
			14'd9460: ff_rdata <= 8'h99;
			14'd9461: ff_rdata <= 8'hF9;
			14'd9462: ff_rdata <= 8'h32;
			14'd9463: ff_rdata <= 8'h97;
			14'd9464: ff_rdata <= 8'hF9;
			14'd9465: ff_rdata <= 8'h32;
			14'd9466: ff_rdata <= 8'h83;
			14'd9467: ff_rdata <= 8'hF9;
			14'd9468: ff_rdata <= 8'h32;
			14'd9469: ff_rdata <= 8'h7F;
			14'd9470: ff_rdata <= 8'hF9;
			14'd9471: ff_rdata <= 8'h32;
			14'd9472: ff_rdata <= 8'h80;
			14'd9473: ff_rdata <= 8'hF9;
			14'd9474: ff_rdata <= 8'h32;
			14'd9475: ff_rdata <= 8'h81;
			14'd9476: ff_rdata <= 8'hF9;
			14'd9477: ff_rdata <= 8'h32;
			14'd9478: ff_rdata <= 8'h82;
			14'd9479: ff_rdata <= 8'hF9;
			14'd9480: ff_rdata <= 8'h6F;
			14'd9481: ff_rdata <= 8'h67;
			14'd9482: ff_rdata <= 8'h22;
			14'd9483: ff_rdata <= 8'h95;
			14'd9484: ff_rdata <= 8'hF9;
			14'd9485: ff_rdata <= 8'h3A;
			14'd9486: ff_rdata <= 8'h91;
			14'd9487: ff_rdata <= 8'hF9;
			14'd9488: ff_rdata <= 8'h47;
			14'd9489: ff_rdata <= 8'h2A;
			14'd9490: ff_rdata <= 8'h7D;
			14'd9491: ff_rdata <= 8'hF9;
			14'd9492: ff_rdata <= 8'h11;
			14'd9493: ff_rdata <= 8'h48;
			14'd9494: ff_rdata <= 8'h00;
			14'd9495: ff_rdata <= 8'h19;
			14'd9496: ff_rdata <= 8'hEB;
			14'd9497: ff_rdata <= 8'hC5;
			14'd9498: ff_rdata <= 8'hD5;
			14'd9499: ff_rdata <= 8'h3A;
			14'd9500: ff_rdata <= 8'h91;
			14'd9501: ff_rdata <= 8'hF9;
			14'd9502: ff_rdata <= 8'h90;
			14'd9503: ff_rdata <= 8'h32;
			14'd9504: ff_rdata <= 8'h9A;
			14'd9505: ff_rdata <= 8'hF9;
			14'd9506: ff_rdata <= 8'h21;
			14'd9507: ff_rdata <= 8'h94;
			14'd9508: ff_rdata <= 8'hF9;
			14'd9509: ff_rdata <= 8'h46;
			14'd9510: ff_rdata <= 8'hCD;
			14'd9511: ff_rdata <= 8'h30;
			14'd9512: ff_rdata <= 8'h67;
			14'd9513: ff_rdata <= 8'hD1;
			14'd9514: ff_rdata <= 8'hC1;
			14'd9515: ff_rdata <= 8'h3A;
			14'd9516: ff_rdata <= 8'h94;
			14'd9517: ff_rdata <= 8'hF9;
			14'd9518: ff_rdata <= 8'h3C;
			14'd9519: ff_rdata <= 8'h6F;
			14'd9520: ff_rdata <= 8'h26;
			14'd9521: ff_rdata <= 8'h00;
			14'd9522: ff_rdata <= 8'h19;
			14'd9523: ff_rdata <= 8'hEB;
			14'd9524: ff_rdata <= 8'h10;
			14'd9525: ff_rdata <= 8'hE3;
			14'd9526: ff_rdata <= 8'h3A;
			14'd9527: ff_rdata <= 8'h92;
			14'd9528: ff_rdata <= 8'hF9;
			14'd9529: ff_rdata <= 8'hB7;
			14'd9530: ff_rdata <= 8'h28;
			14'd9531: ff_rdata <= 8'h15;
			14'd9532: ff_rdata <= 8'h47;
			14'd9533: ff_rdata <= 8'hC5;
			14'd9534: ff_rdata <= 8'h78;
			14'd9535: ff_rdata <= 8'h3D;
			14'd9536: ff_rdata <= 8'h2E;
			14'd9537: ff_rdata <= 8'h00;
			14'd9538: ff_rdata <= 8'hCD;
			14'd9539: ff_rdata <= 8'hE7;
			14'd9540: ff_rdata <= 8'h67;
			14'd9541: ff_rdata <= 8'hEB;
			14'd9542: ff_rdata <= 8'h21;
			14'd9543: ff_rdata <= 8'h66;
			14'd9544: ff_rdata <= 8'h65;
			14'd9545: ff_rdata <= 8'h01;
			14'd9546: ff_rdata <= 8'h27;
			14'd9547: ff_rdata <= 8'h00;
			14'd9548: ff_rdata <= 8'hED;
			14'd9549: ff_rdata <= 8'hB0;
			14'd9550: ff_rdata <= 8'hC1;
			14'd9551: ff_rdata <= 8'h10;
			14'd9552: ff_rdata <= 8'hEC;
			14'd9553: ff_rdata <= 8'hAF;
			14'd9554: ff_rdata <= 8'h32;
			14'd9555: ff_rdata <= 8'h3F;
			14'd9556: ff_rdata <= 8'hFB;
			14'd9557: ff_rdata <= 8'hC9;
			14'd9558: ff_rdata <= 8'h3A;
			14'd9559: ff_rdata <= 8'h8E;
			14'd9560: ff_rdata <= 8'hF9;
			14'd9561: ff_rdata <= 8'hE6;
			14'd9562: ff_rdata <= 8'h01;
			14'd9563: ff_rdata <= 8'hC8;
			14'd9564: ff_rdata <= 8'h3A;
			14'd9565: ff_rdata <= 8'h70;
			14'd9566: ff_rdata <= 8'h65;
			14'd9567: ff_rdata <= 8'h5F;
			14'd9568: ff_rdata <= 8'h3E;
			14'd9569: ff_rdata <= 8'h1F;
			14'd9570: ff_rdata <= 8'hCD;
			14'd9571: ff_rdata <= 8'h2F;
			14'd9572: ff_rdata <= 8'h63;
			14'd9573: ff_rdata <= 8'hC9;
			14'd9574: ff_rdata <= 8'h00;
			14'd9575: ff_rdata <= 8'h00;
			14'd9576: ff_rdata <= 8'h00;
			14'd9577: ff_rdata <= 8'h00;
			14'd9578: ff_rdata <= 8'h00;
			14'd9579: ff_rdata <= 8'h00;
			14'd9580: ff_rdata <= 8'h00;
			14'd9581: ff_rdata <= 8'h00;
			14'd9582: ff_rdata <= 8'h00;
			14'd9583: ff_rdata <= 8'h00;
			14'd9584: ff_rdata <= 8'h0E;
			14'd9585: ff_rdata <= 8'h00;
			14'd9586: ff_rdata <= 8'h00;
			14'd9587: ff_rdata <= 8'h00;
			14'd9588: ff_rdata <= 8'h00;
			14'd9589: ff_rdata <= 8'h04;
			14'd9590: ff_rdata <= 8'h04;
			14'd9591: ff_rdata <= 8'h78;
			14'd9592: ff_rdata <= 8'h08;
			14'd9593: ff_rdata <= 8'h00;
			14'd9594: ff_rdata <= 8'h00;
			14'd9595: ff_rdata <= 8'h00;
			14'd9596: ff_rdata <= 8'h00;
			14'd9597: ff_rdata <= 8'h00;
			14'd9598: ff_rdata <= 8'h00;
			14'd9599: ff_rdata <= 8'h00;
			14'd9600: ff_rdata <= 8'h00;
			14'd9601: ff_rdata <= 8'h00;
			14'd9602: ff_rdata <= 8'h00;
			14'd9603: ff_rdata <= 8'h00;
			14'd9604: ff_rdata <= 8'h00;
			14'd9605: ff_rdata <= 8'h00;
			14'd9606: ff_rdata <= 8'h00;
			14'd9607: ff_rdata <= 8'h00;
			14'd9608: ff_rdata <= 8'h00;
			14'd9609: ff_rdata <= 8'h00;
			14'd9610: ff_rdata <= 8'h00;
			14'd9611: ff_rdata <= 8'h00;
			14'd9612: ff_rdata <= 8'h08;
			14'd9613: ff_rdata <= 8'hCD;
			14'd9614: ff_rdata <= 8'hEE;
			14'd9615: ff_rdata <= 8'h64;
			14'd9616: ff_rdata <= 8'hCD;
			14'd9617: ff_rdata <= 8'h56;
			14'd9618: ff_rdata <= 8'h65;
			14'd9619: ff_rdata <= 8'h3A;
			14'd9620: ff_rdata <= 8'h92;
			14'd9621: ff_rdata <= 8'hF9;
			14'd9622: ff_rdata <= 8'hCD;
			14'd9623: ff_rdata <= 8'h9A;
			14'd9624: ff_rdata <= 8'h65;
			14'd9625: ff_rdata <= 8'hC9;
			14'd9626: ff_rdata <= 8'h3D;
			14'd9627: ff_rdata <= 8'hF8;
			14'd9628: ff_rdata <= 8'h32;
			14'd9629: ff_rdata <= 8'h9A;
			14'd9630: ff_rdata <= 8'hF9;
			14'd9631: ff_rdata <= 8'hF5;
			14'd9632: ff_rdata <= 8'hCD;
			14'd9633: ff_rdata <= 8'h77;
			14'd9634: ff_rdata <= 8'h61;
			14'd9635: ff_rdata <= 8'hF1;
			14'd9636: ff_rdata <= 8'h18;
			14'd9637: ff_rdata <= 8'hF4;
			14'd9638: ff_rdata <= 8'hCD;
			14'd9639: ff_rdata <= 8'hD3;
			14'd9640: ff_rdata <= 8'h67;
			14'd9641: ff_rdata <= 8'hCD;
			14'd9642: ff_rdata <= 8'h34;
			14'd9643: ff_rdata <= 8'h68;
			14'd9644: ff_rdata <= 8'h41;
			14'd9645: ff_rdata <= 8'h4A;
			14'd9646: ff_rdata <= 8'h53;
			14'd9647: ff_rdata <= 8'h78;
			14'd9648: ff_rdata <= 8'hB1;
			14'd9649: ff_rdata <= 8'h28;
			14'd9650: ff_rdata <= 8'h06;
			14'd9651: ff_rdata <= 8'h7A;
			14'd9652: ff_rdata <= 8'hB7;
			14'd9653: ff_rdata <= 8'h28;
			14'd9654: ff_rdata <= 8'h02;
			14'd9655: ff_rdata <= 8'hC5;
			14'd9656: ff_rdata <= 8'hD5;
			14'd9657: ff_rdata <= 8'hF1;
			14'd9658: ff_rdata <= 8'h32;
			14'd9659: ff_rdata <= 8'h3B;
			14'd9660: ff_rdata <= 8'hFB;
			14'd9661: ff_rdata <= 8'hE1;
			14'd9662: ff_rdata <= 8'h7C;
			14'd9663: ff_rdata <= 8'hB5;
			14'd9664: ff_rdata <= 8'hCA;
			14'd9665: ff_rdata <= 8'h15;
			14'd9666: ff_rdata <= 8'h59;
			14'd9667: ff_rdata <= 8'h22;
			14'd9668: ff_rdata <= 8'h3C;
			14'd9669: ff_rdata <= 8'hFB;
			14'd9670: ff_rdata <= 8'hCD;
			14'd9671: ff_rdata <= 8'h1A;
			14'd9672: ff_rdata <= 8'h66;
			14'd9673: ff_rdata <= 8'h28;
			14'd9674: ff_rdata <= 8'hEE;
			14'd9675: ff_rdata <= 8'h2A;
			14'd9676: ff_rdata <= 8'h56;
			14'd9677: ff_rdata <= 8'hF9;
			14'd9678: ff_rdata <= 8'hFE;
			14'd9679: ff_rdata <= 8'h41;
			14'd9680: ff_rdata <= 8'h38;
			14'd9681: ff_rdata <= 8'h04;
			14'd9682: ff_rdata <= 8'hFE;
			14'd9683: ff_rdata <= 8'h48;
			14'd9684: ff_rdata <= 8'h38;
			14'd9685: ff_rdata <= 8'h10;
			14'd9686: ff_rdata <= 8'h87;
			14'd9687: ff_rdata <= 8'h4F;
			14'd9688: ff_rdata <= 8'h7E;
			14'd9689: ff_rdata <= 8'h87;
			14'd9690: ff_rdata <= 8'hCC;
			14'd9691: ff_rdata <= 8'h70;
			14'd9692: ff_rdata <= 8'h67;
			14'd9693: ff_rdata <= 8'hB9;
			14'd9694: ff_rdata <= 8'h28;
			14'd9695: ff_rdata <= 8'h05;
			14'd9696: ff_rdata <= 8'h23;
			14'd9697: ff_rdata <= 8'h23;
			14'd9698: ff_rdata <= 8'h23;
			14'd9699: ff_rdata <= 8'h18;
			14'd9700: ff_rdata <= 8'hF3;
			14'd9701: ff_rdata <= 8'h7E;
			14'd9702: ff_rdata <= 8'h01;
			14'd9703: ff_rdata <= 8'hC6;
			14'd9704: ff_rdata <= 8'h65;
			14'd9705: ff_rdata <= 8'hC5;
			14'd9706: ff_rdata <= 8'h4F;
			14'd9707: ff_rdata <= 8'h87;
			14'd9708: ff_rdata <= 8'h30;
			14'd9709: ff_rdata <= 8'h20;
			14'd9710: ff_rdata <= 8'hB7;
			14'd9711: ff_rdata <= 8'h1F;
			14'd9712: ff_rdata <= 8'h4F;
			14'd9713: ff_rdata <= 8'hC5;
			14'd9714: ff_rdata <= 8'hE5;
			14'd9715: ff_rdata <= 8'hCD;
			14'd9716: ff_rdata <= 8'h1A;
			14'd9717: ff_rdata <= 8'h66;
			14'd9718: ff_rdata <= 8'h11;
			14'd9719: ff_rdata <= 8'h01;
			14'd9720: ff_rdata <= 8'h00;
			14'd9721: ff_rdata <= 8'hCA;
			14'd9722: ff_rdata <= 8'h0B;
			14'd9723: ff_rdata <= 8'h66;
			14'd9724: ff_rdata <= 8'hCD;
			14'd9725: ff_rdata <= 8'hAE;
			14'd9726: ff_rdata <= 8'h68;
			14'd9727: ff_rdata <= 8'hD2;
			14'd9728: ff_rdata <= 8'h08;
			14'd9729: ff_rdata <= 8'h66;
			14'd9730: ff_rdata <= 8'hCD;
			14'd9731: ff_rdata <= 8'h51;
			14'd9732: ff_rdata <= 8'h66;
			14'd9733: ff_rdata <= 8'h37;
			14'd9734: ff_rdata <= 8'h18;
			14'd9735: ff_rdata <= 8'h04;
			14'd9736: ff_rdata <= 8'hCD;
			14'd9737: ff_rdata <= 8'h40;
			14'd9738: ff_rdata <= 8'h66;
			14'd9739: ff_rdata <= 8'hB7;
			14'd9740: ff_rdata <= 8'hE1;
			14'd9741: ff_rdata <= 8'hC1;
			14'd9742: ff_rdata <= 8'h23;
			14'd9743: ff_rdata <= 8'h7E;
			14'd9744: ff_rdata <= 8'h23;
			14'd9745: ff_rdata <= 8'h66;
			14'd9746: ff_rdata <= 8'h6F;
			14'd9747: ff_rdata <= 8'hE9;
			14'd9748: ff_rdata <= 8'hCD;
			14'd9749: ff_rdata <= 8'h1A;
			14'd9750: ff_rdata <= 8'h66;
			14'd9751: ff_rdata <= 8'h28;
			14'd9752: ff_rdata <= 8'hC1;
			14'd9753: ff_rdata <= 8'hC9;
			14'd9754: ff_rdata <= 8'hE5;
			14'd9755: ff_rdata <= 8'h21;
			14'd9756: ff_rdata <= 8'h3B;
			14'd9757: ff_rdata <= 8'hFB;
			14'd9758: ff_rdata <= 8'h7E;
			14'd9759: ff_rdata <= 8'hB7;
			14'd9760: ff_rdata <= 8'h28;
			14'd9761: ff_rdata <= 8'h2A;
			14'd9762: ff_rdata <= 8'h35;
			14'd9763: ff_rdata <= 8'h2A;
			14'd9764: ff_rdata <= 8'h3C;
			14'd9765: ff_rdata <= 8'hFB;
			14'd9766: ff_rdata <= 8'h7E;
			14'd9767: ff_rdata <= 8'h23;
			14'd9768: ff_rdata <= 8'h22;
			14'd9769: ff_rdata <= 8'h3C;
			14'd9770: ff_rdata <= 8'hFB;
			14'd9771: ff_rdata <= 8'hFE;
			14'd9772: ff_rdata <= 8'h20;
			14'd9773: ff_rdata <= 8'h28;
			14'd9774: ff_rdata <= 8'hEC;
			14'd9775: ff_rdata <= 8'hE1;
			14'd9776: ff_rdata <= 8'hCD;
			14'd9777: ff_rdata <= 8'h37;
			14'd9778: ff_rdata <= 8'h66;
			14'd9779: ff_rdata <= 8'h37;
			14'd9780: ff_rdata <= 8'h8F;
			14'd9781: ff_rdata <= 8'h1F;
			14'd9782: ff_rdata <= 8'hC9;
			14'd9783: ff_rdata <= 8'hFE;
			14'd9784: ff_rdata <= 8'h61;
			14'd9785: ff_rdata <= 8'hD8;
			14'd9786: ff_rdata <= 8'hFE;
			14'd9787: ff_rdata <= 8'h7B;
			14'd9788: ff_rdata <= 8'hD0;
			14'd9789: ff_rdata <= 8'hD6;
			14'd9790: ff_rdata <= 8'h20;
			14'd9791: ff_rdata <= 8'hC9;
			14'd9792: ff_rdata <= 8'hE5;
			14'd9793: ff_rdata <= 8'h21;
			14'd9794: ff_rdata <= 8'h3B;
			14'd9795: ff_rdata <= 8'hFB;
			14'd9796: ff_rdata <= 8'h34;
			14'd9797: ff_rdata <= 8'h2A;
			14'd9798: ff_rdata <= 8'h3C;
			14'd9799: ff_rdata <= 8'hFB;
			14'd9800: ff_rdata <= 8'h2B;
			14'd9801: ff_rdata <= 8'h22;
			14'd9802: ff_rdata <= 8'h3C;
			14'd9803: ff_rdata <= 8'hFB;
			14'd9804: ff_rdata <= 8'hE1;
			14'd9805: ff_rdata <= 8'hC9;
			14'd9806: ff_rdata <= 8'hCD;
			14'd9807: ff_rdata <= 8'h14;
			14'd9808: ff_rdata <= 8'h66;
			14'd9809: ff_rdata <= 8'hFE;
			14'd9810: ff_rdata <= 8'h3D;
			14'd9811: ff_rdata <= 8'hCA;
			14'd9812: ff_rdata <= 8'hD3;
			14'd9813: ff_rdata <= 8'h66;
			14'd9814: ff_rdata <= 8'hFE;
			14'd9815: ff_rdata <= 8'h2B;
			14'd9816: ff_rdata <= 8'h28;
			14'd9817: ff_rdata <= 8'hF4;
			14'd9818: ff_rdata <= 8'hFE;
			14'd9819: ff_rdata <= 8'h2D;
			14'd9820: ff_rdata <= 8'h20;
			14'd9821: ff_rdata <= 8'h06;
			14'd9822: ff_rdata <= 8'h11;
			14'd9823: ff_rdata <= 8'hF2;
			14'd9824: ff_rdata <= 8'h66;
			14'd9825: ff_rdata <= 8'hD5;
			14'd9826: ff_rdata <= 8'h18;
			14'd9827: ff_rdata <= 8'hEA;
			14'd9828: ff_rdata <= 8'h11;
			14'd9829: ff_rdata <= 8'h00;
			14'd9830: ff_rdata <= 8'h00;
			14'd9831: ff_rdata <= 8'hFE;
			14'd9832: ff_rdata <= 8'h2C;
			14'd9833: ff_rdata <= 8'h28;
			14'd9834: ff_rdata <= 8'hD5;
			14'd9835: ff_rdata <= 8'hFE;
			14'd9836: ff_rdata <= 8'h3B;
			14'd9837: ff_rdata <= 8'hC8;
			14'd9838: ff_rdata <= 8'hFE;
			14'd9839: ff_rdata <= 8'h3A;
			14'd9840: ff_rdata <= 8'h30;
			14'd9841: ff_rdata <= 8'hCE;
			14'd9842: ff_rdata <= 8'hFE;
			14'd9843: ff_rdata <= 8'h30;
			14'd9844: ff_rdata <= 8'h38;
			14'd9845: ff_rdata <= 8'hCA;
			14'd9846: ff_rdata <= 8'h21;
			14'd9847: ff_rdata <= 8'h00;
			14'd9848: ff_rdata <= 8'h00;
			14'd9849: ff_rdata <= 8'h06;
			14'd9850: ff_rdata <= 8'h0A;
			14'd9851: ff_rdata <= 8'h19;
			14'd9852: ff_rdata <= 8'h38;
			14'd9853: ff_rdata <= 8'h4E;
			14'd9854: ff_rdata <= 8'h10;
			14'd9855: ff_rdata <= 8'hFB;
			14'd9856: ff_rdata <= 8'hD6;
			14'd9857: ff_rdata <= 8'h30;
			14'd9858: ff_rdata <= 8'h5F;
			14'd9859: ff_rdata <= 8'h16;
			14'd9860: ff_rdata <= 8'h00;
			14'd9861: ff_rdata <= 8'h19;
			14'd9862: ff_rdata <= 8'h38;
			14'd9863: ff_rdata <= 8'h44;
			14'd9864: ff_rdata <= 8'hEB;
			14'd9865: ff_rdata <= 8'hCD;
			14'd9866: ff_rdata <= 8'h1A;
			14'd9867: ff_rdata <= 8'h66;
			14'd9868: ff_rdata <= 8'h20;
			14'd9869: ff_rdata <= 8'hD9;
			14'd9870: ff_rdata <= 8'hC9;
			14'd9871: ff_rdata <= 8'hFE;
			14'd9872: ff_rdata <= 8'h41;
			14'd9873: ff_rdata <= 8'hD8;
			14'd9874: ff_rdata <= 8'hFE;
			14'd9875: ff_rdata <= 8'h5B;
			14'd9876: ff_rdata <= 8'h3F;
			14'd9877: ff_rdata <= 8'hC9;
			14'd9878: ff_rdata <= 8'hFE;
			14'd9879: ff_rdata <= 8'h25;
			14'd9880: ff_rdata <= 8'hC8;
			14'd9881: ff_rdata <= 8'hFE;
			14'd9882: ff_rdata <= 8'h21;
			14'd9883: ff_rdata <= 8'hC8;
			14'd9884: ff_rdata <= 8'hFE;
			14'd9885: ff_rdata <= 8'h23;
			14'd9886: ff_rdata <= 8'hC8;
			14'd9887: ff_rdata <= 8'hFE;
			14'd9888: ff_rdata <= 8'h24;
			14'd9889: ff_rdata <= 8'hC8;
			14'd9890: ff_rdata <= 8'h37;
			14'd9891: ff_rdata <= 8'hC9;
			14'd9892: ff_rdata <= 8'hCD;
			14'd9893: ff_rdata <= 8'h14;
			14'd9894: ff_rdata <= 8'h66;
			14'd9895: ff_rdata <= 8'h11;
			14'd9896: ff_rdata <= 8'h5E;
			14'd9897: ff_rdata <= 8'hF5;
			14'd9898: ff_rdata <= 8'hD5;
			14'd9899: ff_rdata <= 8'h06;
			14'd9900: ff_rdata <= 8'h28;
			14'd9901: ff_rdata <= 8'hCD;
			14'd9902: ff_rdata <= 8'h8F;
			14'd9903: ff_rdata <= 8'h66;
			14'd9904: ff_rdata <= 8'h38;
			14'd9905: ff_rdata <= 8'h1A;
			14'd9906: ff_rdata <= 8'h12;
			14'd9907: ff_rdata <= 8'h13;
			14'd9908: ff_rdata <= 8'hCD;
			14'd9909: ff_rdata <= 8'h96;
			14'd9910: ff_rdata <= 8'h66;
			14'd9911: ff_rdata <= 8'h38;
			14'd9912: ff_rdata <= 8'h0A;
			14'd9913: ff_rdata <= 8'hCD;
			14'd9914: ff_rdata <= 8'h14;
			14'd9915: ff_rdata <= 8'h66;
			14'd9916: ff_rdata <= 8'hFE;
			14'd9917: ff_rdata <= 8'h3B;
			14'd9918: ff_rdata <= 8'h20;
			14'd9919: ff_rdata <= 8'h0A;
			14'd9920: ff_rdata <= 8'h12;
			14'd9921: ff_rdata <= 8'h18;
			14'd9922: ff_rdata <= 8'h0C;
			14'd9923: ff_rdata <= 8'hFE;
			14'd9924: ff_rdata <= 8'h3B;
			14'd9925: ff_rdata <= 8'h28;
			14'd9926: ff_rdata <= 8'h08;
			14'd9927: ff_rdata <= 8'hCD;
			14'd9928: ff_rdata <= 8'h14;
			14'd9929: ff_rdata <= 8'h66;
			14'd9930: ff_rdata <= 8'h10;
			14'd9931: ff_rdata <= 8'hE6;
			14'd9932: ff_rdata <= 8'hCD;
			14'd9933: ff_rdata <= 8'h70;
			14'd9934: ff_rdata <= 8'h67;
			14'd9935: ff_rdata <= 8'hE1;
			14'd9936: ff_rdata <= 8'hC3;
			14'd9937: ff_rdata <= 8'h8F;
			14'd9938: ff_rdata <= 8'h67;
			14'd9939: ff_rdata <= 8'hCD;
			14'd9940: ff_rdata <= 8'hA4;
			14'd9941: ff_rdata <= 8'h66;
			14'd9942: ff_rdata <= 8'hCD;
			14'd9943: ff_rdata <= 8'hDE;
			14'd9944: ff_rdata <= 8'hF5;
			14'd9945: ff_rdata <= 8'hEB;
			14'd9946: ff_rdata <= 8'hC9;
			14'd9947: ff_rdata <= 8'hCD;
			14'd9948: ff_rdata <= 8'hA4;
			14'd9949: ff_rdata <= 8'h66;
			14'd9950: ff_rdata <= 8'h3A;
			14'd9951: ff_rdata <= 8'h3B;
			14'd9952: ff_rdata <= 8'hFB;
			14'd9953: ff_rdata <= 8'hB7;
			14'd9954: ff_rdata <= 8'hC2;
			14'd9955: ff_rdata <= 8'h70;
			14'd9956: ff_rdata <= 8'h67;
			14'd9957: ff_rdata <= 8'h2A;
			14'd9958: ff_rdata <= 8'h3C;
			14'd9959: ff_rdata <= 8'hFB;
			14'd9960: ff_rdata <= 8'hE3;
			14'd9961: ff_rdata <= 8'hF5;
			14'd9962: ff_rdata <= 8'h0E;
			14'd9963: ff_rdata <= 8'h02;
			14'd9964: ff_rdata <= 8'hCD;
			14'd9965: ff_rdata <= 8'h94;
			14'd9966: ff_rdata <= 8'h68;
			14'd9967: ff_rdata <= 8'hC3;
			14'd9968: ff_rdata <= 8'hA6;
			14'd9969: ff_rdata <= 8'h65;
			14'd9970: ff_rdata <= 8'hAF;
			14'd9971: ff_rdata <= 8'h93;
			14'd9972: ff_rdata <= 8'h5F;
			14'd9973: ff_rdata <= 8'h9A;
			14'd9974: ff_rdata <= 8'h93;
			14'd9975: ff_rdata <= 8'h57;
			14'd9976: ff_rdata <= 8'hC9;
			14'd9977: ff_rdata <= 8'hCD;
			14'd9978: ff_rdata <= 8'h50;
			14'd9979: ff_rdata <= 8'h67;
			14'd9980: ff_rdata <= 8'h78;
			14'd9981: ff_rdata <= 8'h3C;
			14'd9982: ff_rdata <= 8'h23;
			14'd9983: ff_rdata <= 8'hA6;
			14'd9984: ff_rdata <= 8'hB9;
			14'd9985: ff_rdata <= 8'hC8;
			14'd9986: ff_rdata <= 8'h2B;
			14'd9987: ff_rdata <= 8'h2B;
			14'd9988: ff_rdata <= 8'h2B;
			14'd9989: ff_rdata <= 8'h77;
			14'd9990: ff_rdata <= 8'h23;
			14'd9991: ff_rdata <= 8'h23;
			14'd9992: ff_rdata <= 8'h23;
			14'd9993: ff_rdata <= 8'h23;
			14'd9994: ff_rdata <= 8'h4F;
			14'd9995: ff_rdata <= 8'h7E;
			14'd9996: ff_rdata <= 8'h23;
			14'd9997: ff_rdata <= 8'h66;
			14'd9998: ff_rdata <= 8'h6F;
			14'd9999: ff_rdata <= 8'h06;
			14'd10000: ff_rdata <= 8'h00;
			14'd10001: ff_rdata <= 8'h09;
			14'd10002: ff_rdata <= 8'h73;
			14'd10003: ff_rdata <= 8'hC9;
			14'd10004: ff_rdata <= 8'hCD;
			14'd10005: ff_rdata <= 8'h50;
			14'd10006: ff_rdata <= 8'h67;
			14'd10007: ff_rdata <= 8'h79;
			14'd10008: ff_rdata <= 8'hB8;
			14'd10009: ff_rdata <= 8'hC8;
			14'd10010: ff_rdata <= 8'h23;
			14'd10011: ff_rdata <= 8'h3C;
			14'd10012: ff_rdata <= 8'hA6;
			14'd10013: ff_rdata <= 8'h2B;
			14'd10014: ff_rdata <= 8'h2B;
			14'd10015: ff_rdata <= 8'h77;
			14'd10016: ff_rdata <= 8'h23;
			14'd10017: ff_rdata <= 8'h23;
			14'd10018: ff_rdata <= 8'h23;
			14'd10019: ff_rdata <= 8'h4F;
			14'd10020: ff_rdata <= 8'h7E;
			14'd10021: ff_rdata <= 8'h23;
			14'd10022: ff_rdata <= 8'h66;
			14'd10023: ff_rdata <= 8'h6F;
			14'd10024: ff_rdata <= 8'h06;
			14'd10025: ff_rdata <= 8'h00;
			14'd10026: ff_rdata <= 8'h09;
			14'd10027: ff_rdata <= 8'h7E;
			14'd10028: ff_rdata <= 8'h37;
			14'd10029: ff_rdata <= 8'h8F;
			14'd10030: ff_rdata <= 8'h1F;
			14'd10031: ff_rdata <= 8'hC9;
			14'd10032: ff_rdata <= 8'hC5;
			14'd10033: ff_rdata <= 8'hCD;
			14'd10034: ff_rdata <= 8'h58;
			14'd10035: ff_rdata <= 8'h67;
			14'd10036: ff_rdata <= 8'h70;
			14'd10037: ff_rdata <= 8'h23;
			14'd10038: ff_rdata <= 8'h70;
			14'd10039: ff_rdata <= 8'h23;
			14'd10040: ff_rdata <= 8'h70;
			14'd10041: ff_rdata <= 8'h23;
			14'd10042: ff_rdata <= 8'hF1;
			14'd10043: ff_rdata <= 8'h77;
			14'd10044: ff_rdata <= 8'h23;
			14'd10045: ff_rdata <= 8'h73;
			14'd10046: ff_rdata <= 8'h23;
			14'd10047: ff_rdata <= 8'h72;
			14'd10048: ff_rdata <= 8'hC9;
			14'd10049: ff_rdata <= 8'hCD;
			14'd10050: ff_rdata <= 8'h50;
			14'd10051: ff_rdata <= 8'h67;
			14'd10052: ff_rdata <= 8'h78;
			14'd10053: ff_rdata <= 8'h3C;
			14'd10054: ff_rdata <= 8'h23;
			14'd10055: ff_rdata <= 8'hA6;
			14'd10056: ff_rdata <= 8'h47;
			14'd10057: ff_rdata <= 8'h79;
			14'd10058: ff_rdata <= 8'h90;
			14'd10059: ff_rdata <= 8'hA6;
			14'd10060: ff_rdata <= 8'h6F;
			14'd10061: ff_rdata <= 8'h26;
			14'd10062: ff_rdata <= 8'h00;
			14'd10063: ff_rdata <= 8'hC9;
			14'd10064: ff_rdata <= 8'hCD;
			14'd10065: ff_rdata <= 8'h58;
			14'd10066: ff_rdata <= 8'h67;
			14'd10067: ff_rdata <= 8'h46;
			14'd10068: ff_rdata <= 8'h23;
			14'd10069: ff_rdata <= 8'h4E;
			14'd10070: ff_rdata <= 8'h23;
			14'd10071: ff_rdata <= 8'hC9;
			14'd10072: ff_rdata <= 8'h2A;
			14'd10073: ff_rdata <= 8'h9B;
			14'd10074: ff_rdata <= 8'hF9;
			14'd10075: ff_rdata <= 8'h87;
			14'd10076: ff_rdata <= 8'h47;
			14'd10077: ff_rdata <= 8'h87;
			14'd10078: ff_rdata <= 8'h80;
			14'd10079: ff_rdata <= 8'h4F;
			14'd10080: ff_rdata <= 8'h06;
			14'd10081: ff_rdata <= 8'h00;
			14'd10082: ff_rdata <= 8'h09;
			14'd10083: ff_rdata <= 8'hC9;
			14'd10084: ff_rdata <= 8'h1E;
			14'd10085: ff_rdata <= 8'h33;
			14'd10086: ff_rdata <= 8'h01;
			14'd10087: ff_rdata <= 8'h1E;
			14'd10088: ff_rdata <= 8'h35;
			14'd10089: ff_rdata <= 8'h01;
			14'd10090: ff_rdata <= 8'h1E;
			14'd10091: ff_rdata <= 8'h38;
			14'd10092: ff_rdata <= 8'h01;
			14'd10093: ff_rdata <= 8'h1E;
			14'd10094: ff_rdata <= 8'h02;
			14'd10095: ff_rdata <= 8'h01;
			14'd10096: ff_rdata <= 8'h1E;
			14'd10097: ff_rdata <= 8'h05;
			14'd10098: ff_rdata <= 8'h01;
			14'd10099: ff_rdata <= 8'h1E;
			14'd10100: ff_rdata <= 8'h0D;
			14'd10101: ff_rdata <= 8'h01;
			14'd10102: ff_rdata <= 8'h1E;
			14'd10103: ff_rdata <= 8'h06;
			14'd10104: ff_rdata <= 8'h01;
			14'd10105: ff_rdata <= 8'h1E;
			14'd10106: ff_rdata <= 8'h07;
			14'd10107: ff_rdata <= 8'hCD;
			14'd10108: ff_rdata <= 8'hC6;
			14'd10109: ff_rdata <= 8'h50;
			14'd10110: ff_rdata <= 8'hD5;
			14'd10111: ff_rdata <= 8'hC4;
			14'd10112: ff_rdata <= 8'h8D;
			14'd10113: ff_rdata <= 8'h65;
			14'd10114: ff_rdata <= 8'hD1;
			14'd10115: ff_rdata <= 8'hDD;
			14'd10116: ff_rdata <= 8'h21;
			14'd10117: ff_rdata <= 8'h6F;
			14'd10118: ff_rdata <= 8'h40;
			14'd10119: ff_rdata <= 8'h18;
			14'd10120: ff_rdata <= 8'h4E;
			14'd10121: ff_rdata <= 8'hDD;
			14'd10122: ff_rdata <= 8'h21;
			14'd10123: ff_rdata <= 8'h90;
			14'd10124: ff_rdata <= 8'h00;
			14'd10125: ff_rdata <= 8'h18;
			14'd10126: ff_rdata <= 8'h48;
			14'd10127: ff_rdata <= 8'hDD;
			14'd10128: ff_rdata <= 8'h21;
			14'd10129: ff_rdata <= 8'h9B;
			14'd10130: ff_rdata <= 8'h4E;
			14'd10131: ff_rdata <= 8'h18;
			14'd10132: ff_rdata <= 8'h42;
			14'd10133: ff_rdata <= 8'hDD;
			14'd10134: ff_rdata <= 8'h21;
			14'd10135: ff_rdata <= 8'h0E;
			14'd10136: ff_rdata <= 8'h6A;
			14'd10137: ff_rdata <= 8'h18;
			14'd10138: ff_rdata <= 8'h3C;
			14'd10139: ff_rdata <= 8'hDD;
			14'd10140: ff_rdata <= 8'h21;
			14'd10141: ff_rdata <= 8'hA4;
			14'd10142: ff_rdata <= 8'h5E;
			14'd10143: ff_rdata <= 8'h18;
			14'd10144: ff_rdata <= 8'h36;
			14'd10145: ff_rdata <= 8'hDD;
			14'd10146: ff_rdata <= 8'h21;
			14'd10147: ff_rdata <= 8'h7A;
			14'd10148: ff_rdata <= 8'h51;
			14'd10149: ff_rdata <= 8'h18;
			14'd10150: ff_rdata <= 8'h30;
			14'd10151: ff_rdata <= 8'h7E;
			14'd10152: ff_rdata <= 8'hE3;
			14'd10153: ff_rdata <= 8'hBE;
			14'd10154: ff_rdata <= 8'hC2;
			14'd10155: ff_rdata <= 8'h6D;
			14'd10156: ff_rdata <= 8'h67;
			14'd10157: ff_rdata <= 8'h23;
			14'd10158: ff_rdata <= 8'hE3;
			14'd10159: ff_rdata <= 8'hDD;
			14'd10160: ff_rdata <= 8'h21;
			14'd10161: ff_rdata <= 8'h66;
			14'd10162: ff_rdata <= 8'h46;
			14'd10163: ff_rdata <= 8'h18;
			14'd10164: ff_rdata <= 8'h22;
			14'd10165: ff_rdata <= 8'hDD;
			14'd10166: ff_rdata <= 8'h21;
			14'd10167: ff_rdata <= 8'h64;
			14'd10168: ff_rdata <= 8'h4C;
			14'd10169: ff_rdata <= 8'h18;
			14'd10170: ff_rdata <= 8'h1C;
			14'd10171: ff_rdata <= 8'hDD;
			14'd10172: ff_rdata <= 8'h21;
			14'd10173: ff_rdata <= 8'h2F;
			14'd10174: ff_rdata <= 8'h54;
			14'd10175: ff_rdata <= 8'h18;
			14'd10176: ff_rdata <= 8'h16;
			14'd10177: ff_rdata <= 8'hDD;
			14'd10178: ff_rdata <= 8'h21;
			14'd10179: ff_rdata <= 8'h1C;
			14'd10180: ff_rdata <= 8'h52;
			14'd10181: ff_rdata <= 8'h18;
			14'd10182: ff_rdata <= 8'h10;
			14'd10183: ff_rdata <= 8'hDD;
			14'd10184: ff_rdata <= 8'h21;
			14'd10185: ff_rdata <= 8'h01;
			14'd10186: ff_rdata <= 8'h46;
			14'd10187: ff_rdata <= 8'h18;
			14'd10188: ff_rdata <= 8'h0A;
			14'd10189: ff_rdata <= 8'hDD;
			14'd10190: ff_rdata <= 8'h21;
			14'd10191: ff_rdata <= 8'h1C;
			14'd10192: ff_rdata <= 8'h6C;
			14'd10193: ff_rdata <= 8'h18;
			14'd10194: ff_rdata <= 8'h04;
			14'd10195: ff_rdata <= 8'hDD;
			14'd10196: ff_rdata <= 8'h21;
			14'd10197: ff_rdata <= 8'hD0;
			14'd10198: ff_rdata <= 8'h67;
			14'd10199: ff_rdata <= 8'hFD;
			14'd10200: ff_rdata <= 8'h2A;
			14'd10201: ff_rdata <= 8'hC0;
			14'd10202: ff_rdata <= 8'hFC;
			14'd10203: ff_rdata <= 8'hCD;
			14'd10204: ff_rdata <= 8'h1C;
			14'd10205: ff_rdata <= 8'h00;
			14'd10206: ff_rdata <= 8'hFB;
			14'd10207: ff_rdata <= 8'hC9;
			14'd10208: ff_rdata <= 8'h2E;
			14'd10209: ff_rdata <= 8'h02;
			14'd10210: ff_rdata <= 8'h18;
			14'd10211: ff_rdata <= 8'h03;
			14'd10212: ff_rdata <= 8'h3A;
			14'd10213: ff_rdata <= 8'h38;
			14'd10214: ff_rdata <= 8'hFB;
			14'd10215: ff_rdata <= 8'h26;
			14'd10216: ff_rdata <= 8'h00;
			14'd10217: ff_rdata <= 8'hD5;
			14'd10218: ff_rdata <= 8'h5F;
			14'd10219: ff_rdata <= 8'h3A;
			14'd10220: ff_rdata <= 8'h91;
			14'd10221: ff_rdata <= 8'hF9;
			14'd10222: ff_rdata <= 8'h93;
			14'd10223: ff_rdata <= 8'hD6;
			14'd10224: ff_rdata <= 8'h04;
			14'd10225: ff_rdata <= 8'h38;
			14'd10226: ff_rdata <= 8'h12;
			14'd10227: ff_rdata <= 8'h7B;
			14'd10228: ff_rdata <= 8'h11;
			14'd10229: ff_rdata <= 8'hC8;
			14'd10230: ff_rdata <= 8'h01;
			14'd10231: ff_rdata <= 8'h19;
			14'd10232: ff_rdata <= 8'hED;
			14'd10233: ff_rdata <= 8'h5B;
			14'd10234: ff_rdata <= 8'h7D;
			14'd10235: ff_rdata <= 8'hF9;
			14'd10236: ff_rdata <= 8'h19;
			14'd10237: ff_rdata <= 8'hB7;
			14'd10238: ff_rdata <= 8'h28;
			14'd10239: ff_rdata <= 8'h25;
			14'd10240: ff_rdata <= 8'h11;
			14'd10241: ff_rdata <= 8'h27;
			14'd10242: ff_rdata <= 8'h00;
			14'd10243: ff_rdata <= 8'h18;
			14'd10244: ff_rdata <= 8'h1C;
			14'd10245: ff_rdata <= 8'h2F;
			14'd10246: ff_rdata <= 8'h08;
			14'd10247: ff_rdata <= 8'h7D;
			14'd10248: ff_rdata <= 8'hB7;
			14'd10249: ff_rdata <= 8'h20;
			14'd10250: ff_rdata <= 8'h0B;
			14'd10251: ff_rdata <= 8'h08;
			14'd10252: ff_rdata <= 8'h21;
			14'd10253: ff_rdata <= 8'hAF;
			14'd10254: ff_rdata <= 8'hF9;
			14'd10255: ff_rdata <= 8'h87;
			14'd10256: ff_rdata <= 8'hCD;
			14'd10257: ff_rdata <= 8'h86;
			14'd10258: ff_rdata <= 8'h54;
			14'd10259: ff_rdata <= 8'hD1;
			14'd10260: ff_rdata <= 8'hAF;
			14'd10261: ff_rdata <= 8'hC9;
			14'd10262: ff_rdata <= 8'h08;
			14'd10263: ff_rdata <= 8'h11;
			14'd10264: ff_rdata <= 8'h41;
			14'd10265: ff_rdata <= 8'hFB;
			14'd10266: ff_rdata <= 8'h19;
			14'd10267: ff_rdata <= 8'hB7;
			14'd10268: ff_rdata <= 8'h28;
			14'd10269: ff_rdata <= 8'h07;
			14'd10270: ff_rdata <= 8'h11;
			14'd10271: ff_rdata <= 8'h25;
			14'd10272: ff_rdata <= 8'h00;
			14'd10273: ff_rdata <= 8'h19;
			14'd10274: ff_rdata <= 8'h3D;
			14'd10275: ff_rdata <= 8'h20;
			14'd10276: ff_rdata <= 8'hFC;
			14'd10277: ff_rdata <= 8'hD1;
			14'd10278: ff_rdata <= 8'hC9;
			14'd10279: ff_rdata <= 8'hC5;
			14'd10280: ff_rdata <= 8'hE3;
			14'd10281: ff_rdata <= 8'hC1;
			14'd10282: ff_rdata <= 8'hCD;
			14'd10283: ff_rdata <= 8'hD4;
			14'd10284: ff_rdata <= 8'h68;
			14'd10285: ff_rdata <= 8'h7E;
			14'd10286: ff_rdata <= 8'h02;
			14'd10287: ff_rdata <= 8'hC8;
			14'd10288: ff_rdata <= 8'h0B;
			14'd10289: ff_rdata <= 8'h2B;
			14'd10290: ff_rdata <= 8'h18;
			14'd10291: ff_rdata <= 8'hF6;
			14'd10292: ff_rdata <= 8'h5E;
			14'd10293: ff_rdata <= 8'h23;
			14'd10294: ff_rdata <= 8'h56;
			14'd10295: ff_rdata <= 8'h23;
			14'd10296: ff_rdata <= 8'h4E;
			14'd10297: ff_rdata <= 8'h23;
			14'd10298: ff_rdata <= 8'h46;
			14'd10299: ff_rdata <= 8'h23;
			14'd10300: ff_rdata <= 8'hC9;
			14'd10301: ff_rdata <= 8'hF3;
			14'd10302: ff_rdata <= 8'h2A;
			14'd10303: ff_rdata <= 8'h95;
			14'd10304: ff_rdata <= 8'hF9;
			14'd10305: ff_rdata <= 8'h7D;
			14'd10306: ff_rdata <= 8'hB4;
			14'd10307: ff_rdata <= 8'hC0;
			14'd10308: ff_rdata <= 8'h21;
			14'd10309: ff_rdata <= 8'h40;
			14'd10310: ff_rdata <= 8'hFB;
			14'd10311: ff_rdata <= 8'hB6;
			14'd10312: ff_rdata <= 8'h28;
			14'd10313: ff_rdata <= 8'h1D;
			14'd10314: ff_rdata <= 8'h35;
			14'd10315: ff_rdata <= 8'h21;
			14'd10316: ff_rdata <= 8'hFF;
			14'd10317: ff_rdata <= 8'hFF;
			14'd10318: ff_rdata <= 8'h22;
			14'd10319: ff_rdata <= 8'h41;
			14'd10320: ff_rdata <= 8'hFB;
			14'd10321: ff_rdata <= 8'h22;
			14'd10322: ff_rdata <= 8'h66;
			14'd10323: ff_rdata <= 8'hFB;
			14'd10324: ff_rdata <= 8'h22;
			14'd10325: ff_rdata <= 8'h8B;
			14'd10326: ff_rdata <= 8'hFB;
			14'd10327: ff_rdata <= 8'h23;
			14'd10328: ff_rdata <= 8'h23;
			14'd10329: ff_rdata <= 8'h22;
			14'd10330: ff_rdata <= 8'hAF;
			14'd10331: ff_rdata <= 8'hF9;
			14'd10332: ff_rdata <= 8'h22;
			14'd10333: ff_rdata <= 8'hB1;
			14'd10334: ff_rdata <= 8'hF9;
			14'd10335: ff_rdata <= 8'h22;
			14'd10336: ff_rdata <= 8'hB3;
			14'd10337: ff_rdata <= 8'hF9;
			14'd10338: ff_rdata <= 8'h3E;
			14'd10339: ff_rdata <= 8'h87;
			14'd10340: ff_rdata <= 8'h32;
			14'd10341: ff_rdata <= 8'h3F;
			14'd10342: ff_rdata <= 8'hFB;
			14'd10343: ff_rdata <= 8'h21;
			14'd10344: ff_rdata <= 8'h97;
			14'd10345: ff_rdata <= 8'hF9;
			14'd10346: ff_rdata <= 8'h7E;
			14'd10347: ff_rdata <= 8'hB7;
			14'd10348: ff_rdata <= 8'hC8;
			14'd10349: ff_rdata <= 8'h35;
			14'd10350: ff_rdata <= 8'h3A;
			14'd10351: ff_rdata <= 8'h92;
			14'd10352: ff_rdata <= 8'hF9;
			14'd10353: ff_rdata <= 8'hB7;
			14'd10354: ff_rdata <= 8'h28;
			14'd10355: ff_rdata <= 8'h14;
			14'd10356: ff_rdata <= 8'h47;
			14'd10357: ff_rdata <= 8'h2A;
			14'd10358: ff_rdata <= 8'h7D;
			14'd10359: ff_rdata <= 8'hF9;
			14'd10360: ff_rdata <= 8'h11;
			14'd10361: ff_rdata <= 8'hC8;
			14'd10362: ff_rdata <= 8'h01;
			14'd10363: ff_rdata <= 8'h19;
			14'd10364: ff_rdata <= 8'h11;
			14'd10365: ff_rdata <= 8'h27;
			14'd10366: ff_rdata <= 8'h00;
			14'd10367: ff_rdata <= 8'h36;
			14'd10368: ff_rdata <= 8'h01;
			14'd10369: ff_rdata <= 8'h23;
			14'd10370: ff_rdata <= 8'h36;
			14'd10371: ff_rdata <= 8'h00;
			14'd10372: ff_rdata <= 8'h2B;
			14'd10373: ff_rdata <= 8'h19;
			14'd10374: ff_rdata <= 8'h10;
			14'd10375: ff_rdata <= 8'hF7;
			14'd10376: ff_rdata <= 8'h2A;
			14'd10377: ff_rdata <= 8'h8F;
			14'd10378: ff_rdata <= 8'hF9;
			14'd10379: ff_rdata <= 8'h22;
			14'd10380: ff_rdata <= 8'h95;
			14'd10381: ff_rdata <= 8'hF9;
			14'd10382: ff_rdata <= 8'h3E;
			14'd10383: ff_rdata <= 8'hFF;
			14'd10384: ff_rdata <= 8'h32;
			14'd10385: ff_rdata <= 8'h26;
			14'd10386: ff_rdata <= 8'hFA;
			14'd10387: ff_rdata <= 8'hC9;
			14'd10388: ff_rdata <= 8'hE5;
			14'd10389: ff_rdata <= 8'h2A;
			14'd10390: ff_rdata <= 8'hC6;
			14'd10391: ff_rdata <= 8'hF6;
			14'd10392: ff_rdata <= 8'h06;
			14'd10393: ff_rdata <= 8'h00;
			14'd10394: ff_rdata <= 8'h09;
			14'd10395: ff_rdata <= 8'h09;
			14'd10396: ff_rdata <= 8'h3E;
			14'd10397: ff_rdata <= 8'hE5;
			14'd10398: ff_rdata <= 8'h3E;
			14'd10399: ff_rdata <= 8'h88;
			14'd10400: ff_rdata <= 8'h95;
			14'd10401: ff_rdata <= 8'h6F;
			14'd10402: ff_rdata <= 8'h3E;
			14'd10403: ff_rdata <= 8'hFF;
			14'd10404: ff_rdata <= 8'h9C;
			14'd10405: ff_rdata <= 8'h67;
			14'd10406: ff_rdata <= 8'h38;
			14'd10407: ff_rdata <= 8'h03;
			14'd10408: ff_rdata <= 8'h39;
			14'd10409: ff_rdata <= 8'hE1;
			14'd10410: ff_rdata <= 8'hD8;
			14'd10411: ff_rdata <= 8'hC3;
			14'd10412: ff_rdata <= 8'h79;
			14'd10413: ff_rdata <= 8'h67;
			14'd10414: ff_rdata <= 8'hFE;
			14'd10415: ff_rdata <= 8'h7B;
			14'd10416: ff_rdata <= 8'hC8;
			14'd10417: ff_rdata <= 8'hFE;
			14'd10418: ff_rdata <= 8'h7D;
			14'd10419: ff_rdata <= 8'hC8;
			14'd10420: ff_rdata <= 8'hFE;
			14'd10421: ff_rdata <= 8'h3E;
			14'd10422: ff_rdata <= 8'hC8;
			14'd10423: ff_rdata <= 8'hFE;
			14'd10424: ff_rdata <= 8'h3C;
			14'd10425: ff_rdata <= 8'hC8;
			14'd10426: ff_rdata <= 8'hFE;
			14'd10427: ff_rdata <= 8'h26;
			14'd10428: ff_rdata <= 8'hC8;
			14'd10429: ff_rdata <= 8'hFE;
			14'd10430: ff_rdata <= 8'h40;
			14'd10431: ff_rdata <= 8'hD8;
			14'd10432: ff_rdata <= 8'hFE;
			14'd10433: ff_rdata <= 8'h5B;
			14'd10434: ff_rdata <= 8'h3F;
			14'd10435: ff_rdata <= 8'hC9;
			14'd10436: ff_rdata <= 8'h3A;
			14'd10437: ff_rdata <= 8'h63;
			14'd10438: ff_rdata <= 8'hF6;
			14'd10439: ff_rdata <= 8'hFE;
			14'd10440: ff_rdata <= 8'h08;
			14'd10441: ff_rdata <= 8'h30;
			14'd10442: ff_rdata <= 8'h05;
			14'd10443: ff_rdata <= 8'hD6;
			14'd10444: ff_rdata <= 8'h03;
			14'd10445: ff_rdata <= 8'hB7;
			14'd10446: ff_rdata <= 8'h37;
			14'd10447: ff_rdata <= 8'hC9;
			14'd10448: ff_rdata <= 8'hD6;
			14'd10449: ff_rdata <= 8'h03;
			14'd10450: ff_rdata <= 8'hB7;
			14'd10451: ff_rdata <= 8'hC9;
			14'd10452: ff_rdata <= 8'h7C;
			14'd10453: ff_rdata <= 8'h92;
			14'd10454: ff_rdata <= 8'hC0;
			14'd10455: ff_rdata <= 8'h7D;
			14'd10456: ff_rdata <= 8'h93;
			14'd10457: ff_rdata <= 8'hC9;
			14'd10458: ff_rdata <= 8'h69;
			14'd10459: ff_rdata <= 8'h60;
			14'd10460: ff_rdata <= 8'hCD;
			14'd10461: ff_rdata <= 8'h42;
			14'd10462: ff_rdata <= 8'h69;
			14'd10463: ff_rdata <= 8'h18;
			14'd10464: ff_rdata <= 8'h12;
			14'd10465: ff_rdata <= 8'h79;
			14'd10466: ff_rdata <= 8'hFE;
			14'd10467: ff_rdata <= 8'h40;
			14'd10468: ff_rdata <= 8'hD0;
			14'd10469: ff_rdata <= 8'hCD;
			14'd10470: ff_rdata <= 8'h0F;
			14'd10471: ff_rdata <= 8'h69;
			14'd10472: ff_rdata <= 8'hDD;
			14'd10473: ff_rdata <= 8'h36;
			14'd10474: ff_rdata <= 8'h07;
			14'd10475: ff_rdata <= 8'h00;
			14'd10476: ff_rdata <= 8'hDD;
			14'd10477: ff_rdata <= 8'h36;
			14'd10478: ff_rdata <= 8'h08;
			14'd10479: ff_rdata <= 8'h00;
			14'd10480: ff_rdata <= 8'hC4;
			14'd10481: ff_rdata <= 8'h38;
			14'd10482: ff_rdata <= 8'h69;
			14'd10483: ff_rdata <= 8'hC5;
			14'd10484: ff_rdata <= 8'hDD;
			14'd10485: ff_rdata <= 8'h7E;
			14'd10486: ff_rdata <= 8'h00;
			14'd10487: ff_rdata <= 8'hC6;
			14'd10488: ff_rdata <= 8'h20;
			14'd10489: ff_rdata <= 8'h4F;
			14'd10490: ff_rdata <= 8'hCD;
			14'd10491: ff_rdata <= 8'hE0;
			14'd10492: ff_rdata <= 8'h6D;
			14'd10493: ff_rdata <= 8'hE6;
			14'd10494: ff_rdata <= 8'h0F;
			14'd10495: ff_rdata <= 8'h47;
			14'd10496: ff_rdata <= 8'hD1;
			14'd10497: ff_rdata <= 8'h7B;
			14'd10498: ff_rdata <= 8'h87;
			14'd10499: ff_rdata <= 8'h87;
			14'd10500: ff_rdata <= 8'h87;
			14'd10501: ff_rdata <= 8'h87;
			14'd10502: ff_rdata <= 8'hB0;
			14'd10503: ff_rdata <= 8'h47;
			14'd10504: ff_rdata <= 8'hCD;
			14'd10505: ff_rdata <= 8'hB5;
			14'd10506: ff_rdata <= 8'h6D;
			14'd10507: ff_rdata <= 8'hCD;
			14'd10508: ff_rdata <= 8'h78;
			14'd10509: ff_rdata <= 8'h6A;
			14'd10510: ff_rdata <= 8'hC9;
			14'd10511: ff_rdata <= 8'hC5;
			14'd10512: ff_rdata <= 8'hE5;
			14'd10513: ff_rdata <= 8'h21;
			14'd10514: ff_rdata <= 8'h28;
			14'd10515: ff_rdata <= 8'h69;
			14'd10516: ff_rdata <= 8'h79;
			14'd10517: ff_rdata <= 8'h01;
			14'd10518: ff_rdata <= 8'h10;
			14'd10519: ff_rdata <= 8'h00;
			14'd10520: ff_rdata <= 8'hED;
			14'd10521: ff_rdata <= 8'hB1;
			14'd10522: ff_rdata <= 8'h28;
			14'd10523: ff_rdata <= 8'h03;
			14'd10524: ff_rdata <= 8'hE1;
			14'd10525: ff_rdata <= 8'hC1;
			14'd10526: ff_rdata <= 8'hC9;
			14'd10527: ff_rdata <= 8'h3E;
			14'd10528: ff_rdata <= 8'h10;
			14'd10529: ff_rdata <= 8'h91;
			14'd10530: ff_rdata <= 8'h3D;
			14'd10531: ff_rdata <= 8'hE1;
			14'd10532: ff_rdata <= 8'hC1;
			14'd10533: ff_rdata <= 8'h4F;
			14'd10534: ff_rdata <= 8'hAF;
			14'd10535: ff_rdata <= 8'hC9;
			14'd10536: ff_rdata <= 8'hFF;
			14'd10537: ff_rdata <= 8'h02;
			14'd10538: ff_rdata <= 8'h0A;
			14'd10539: ff_rdata <= 8'h00;
			14'd10540: ff_rdata <= 8'h03;
			14'd10541: ff_rdata <= 8'h04;
			14'd10542: ff_rdata <= 8'h05;
			14'd10543: ff_rdata <= 8'h06;
			14'd10544: ff_rdata <= 8'h09;
			14'd10545: ff_rdata <= 8'h30;
			14'd10546: ff_rdata <= 8'h18;
			14'd10547: ff_rdata <= 8'h0E;
			14'd10548: ff_rdata <= 8'h10;
			14'd10549: ff_rdata <= 8'h17;
			14'd10550: ff_rdata <= 8'h21;
			14'd10551: ff_rdata <= 8'h0C;
			14'd10552: ff_rdata <= 8'hE5;
			14'd10553: ff_rdata <= 8'h69;
			14'd10554: ff_rdata <= 8'hCD;
			14'd10555: ff_rdata <= 8'h32;
			14'd10556: ff_rdata <= 8'h57;
			14'd10557: ff_rdata <= 8'hCD;
			14'd10558: ff_rdata <= 8'h42;
			14'd10559: ff_rdata <= 8'h69;
			14'd10560: ff_rdata <= 8'hE1;
			14'd10561: ff_rdata <= 8'hC9;
			14'd10562: ff_rdata <= 8'h11;
			14'd10563: ff_rdata <= 8'h08;
			14'd10564: ff_rdata <= 8'h00;
			14'd10565: ff_rdata <= 8'h19;
			14'd10566: ff_rdata <= 8'h5E;
			14'd10567: ff_rdata <= 8'h23;
			14'd10568: ff_rdata <= 8'h56;
			14'd10569: ff_rdata <= 8'h23;
			14'd10570: ff_rdata <= 8'hDD;
			14'd10571: ff_rdata <= 8'h73;
			14'd10572: ff_rdata <= 8'h07;
			14'd10573: ff_rdata <= 8'hDD;
			14'd10574: ff_rdata <= 8'h72;
			14'd10575: ff_rdata <= 8'h08;
			14'd10576: ff_rdata <= 8'hDD;
			14'd10577: ff_rdata <= 8'hE5;
			14'd10578: ff_rdata <= 8'hDD;
			14'd10579: ff_rdata <= 8'h21;
			14'd10580: ff_rdata <= 8'h27;
			14'd10581: ff_rdata <= 8'hFA;
			14'd10582: ff_rdata <= 8'h06;
			14'd10583: ff_rdata <= 8'h09;
			14'd10584: ff_rdata <= 8'hC5;
			14'd10585: ff_rdata <= 8'hDD;
			14'd10586: ff_rdata <= 8'h7E;
			14'd10587: ff_rdata <= 8'h00;
			14'd10588: ff_rdata <= 8'hC6;
			14'd10589: ff_rdata <= 8'h20;
			14'd10590: ff_rdata <= 8'h4F;
			14'd10591: ff_rdata <= 8'hCD;
			14'd10592: ff_rdata <= 8'hE0;
			14'd10593: ff_rdata <= 8'h6D;
			14'd10594: ff_rdata <= 8'h0F;
			14'd10595: ff_rdata <= 8'h0F;
			14'd10596: ff_rdata <= 8'h0F;
			14'd10597: ff_rdata <= 8'h0F;
			14'd10598: ff_rdata <= 8'hE6;
			14'd10599: ff_rdata <= 8'h0F;
			14'd10600: ff_rdata <= 8'h20;
			14'd10601: ff_rdata <= 8'h06;
			14'd10602: ff_rdata <= 8'hDD;
			14'd10603: ff_rdata <= 8'h73;
			14'd10604: ff_rdata <= 8'h07;
			14'd10605: ff_rdata <= 8'hDD;
			14'd10606: ff_rdata <= 8'h72;
			14'd10607: ff_rdata <= 8'h08;
			14'd10608: ff_rdata <= 8'h01;
			14'd10609: ff_rdata <= 8'h10;
			14'd10610: ff_rdata <= 8'h00;
			14'd10611: ff_rdata <= 8'hDD;
			14'd10612: ff_rdata <= 8'h09;
			14'd10613: ff_rdata <= 8'hC1;
			14'd10614: ff_rdata <= 8'h10;
			14'd10615: ff_rdata <= 8'hE0;
			14'd10616: ff_rdata <= 8'hDD;
			14'd10617: ff_rdata <= 8'hE1;
			14'd10618: ff_rdata <= 8'h7E;
			14'd10619: ff_rdata <= 8'h11;
			14'd10620: ff_rdata <= 8'h06;
			14'd10621: ff_rdata <= 8'h00;
			14'd10622: ff_rdata <= 8'h19;
			14'd10623: ff_rdata <= 8'hE6;
			14'd10624: ff_rdata <= 8'h0E;
			14'd10625: ff_rdata <= 8'h0F;
			14'd10626: ff_rdata <= 8'h57;
			14'd10627: ff_rdata <= 8'h46;
			14'd10628: ff_rdata <= 8'h0E;
			14'd10629: ff_rdata <= 8'h00;
			14'd10630: ff_rdata <= 8'hCD;
			14'd10631: ff_rdata <= 8'hB5;
			14'd10632: ff_rdata <= 8'h6D;
			14'd10633: ff_rdata <= 8'h23;
			14'd10634: ff_rdata <= 8'h46;
			14'd10635: ff_rdata <= 8'h0E;
			14'd10636: ff_rdata <= 8'h02;
			14'd10637: ff_rdata <= 8'hCD;
			14'd10638: ff_rdata <= 8'hB5;
			14'd10639: ff_rdata <= 8'h6D;
			14'd10640: ff_rdata <= 8'h23;
			14'd10641: ff_rdata <= 8'h46;
			14'd10642: ff_rdata <= 8'h0E;
			14'd10643: ff_rdata <= 8'h04;
			14'd10644: ff_rdata <= 8'hCD;
			14'd10645: ff_rdata <= 8'hB5;
			14'd10646: ff_rdata <= 8'h6D;
			14'd10647: ff_rdata <= 8'h23;
			14'd10648: ff_rdata <= 8'h46;
			14'd10649: ff_rdata <= 8'h0E;
			14'd10650: ff_rdata <= 8'h06;
			14'd10651: ff_rdata <= 8'hCD;
			14'd10652: ff_rdata <= 8'hB5;
			14'd10653: ff_rdata <= 8'h6D;
			14'd10654: ff_rdata <= 8'h23;
			14'd10655: ff_rdata <= 8'h23;
			14'd10656: ff_rdata <= 8'h23;
			14'd10657: ff_rdata <= 8'h23;
			14'd10658: ff_rdata <= 8'h23;
			14'd10659: ff_rdata <= 8'h46;
			14'd10660: ff_rdata <= 8'h0E;
			14'd10661: ff_rdata <= 8'h01;
			14'd10662: ff_rdata <= 8'hCD;
			14'd10663: ff_rdata <= 8'hB5;
			14'd10664: ff_rdata <= 8'h6D;
			14'd10665: ff_rdata <= 8'h23;
			14'd10666: ff_rdata <= 8'h7E;
			14'd10667: ff_rdata <= 8'hE6;
			14'd10668: ff_rdata <= 8'hC0;
			14'd10669: ff_rdata <= 8'hB2;
			14'd10670: ff_rdata <= 8'h57;
			14'd10671: ff_rdata <= 8'h0E;
			14'd10672: ff_rdata <= 8'h03;
			14'd10673: ff_rdata <= 8'hCD;
			14'd10674: ff_rdata <= 8'hE0;
			14'd10675: ff_rdata <= 8'h6D;
			14'd10676: ff_rdata <= 8'hE6;
			14'd10677: ff_rdata <= 8'h18;
			14'd10678: ff_rdata <= 8'hB2;
			14'd10679: ff_rdata <= 8'h47;
			14'd10680: ff_rdata <= 8'hCD;
			14'd10681: ff_rdata <= 8'hB5;
			14'd10682: ff_rdata <= 8'h6D;
			14'd10683: ff_rdata <= 8'h23;
			14'd10684: ff_rdata <= 8'h46;
			14'd10685: ff_rdata <= 8'h0E;
			14'd10686: ff_rdata <= 8'h05;
			14'd10687: ff_rdata <= 8'hCD;
			14'd10688: ff_rdata <= 8'hB5;
			14'd10689: ff_rdata <= 8'h6D;
			14'd10690: ff_rdata <= 8'h23;
			14'd10691: ff_rdata <= 8'h46;
			14'd10692: ff_rdata <= 8'h0E;
			14'd10693: ff_rdata <= 8'h07;
			14'd10694: ff_rdata <= 8'hCD;
			14'd10695: ff_rdata <= 8'hB5;
			14'd10696: ff_rdata <= 8'h6D;
			14'd10697: ff_rdata <= 8'h0E;
			14'd10698: ff_rdata <= 8'h00;
			14'd10699: ff_rdata <= 8'hC9;
			14'd10700: ff_rdata <= 8'h7B;
			14'd10701: ff_rdata <= 8'h0F;
			14'd10702: ff_rdata <= 8'h0F;
			14'd10703: ff_rdata <= 8'h0F;
			14'd10704: ff_rdata <= 8'hE6;
			14'd10705: ff_rdata <= 8'h07;
			14'd10706: ff_rdata <= 8'hDD;
			14'd10707: ff_rdata <= 8'h77;
			14'd10708: ff_rdata <= 8'h02;
			14'd10709: ff_rdata <= 8'hE5;
			14'd10710: ff_rdata <= 8'hCD;
			14'd10711: ff_rdata <= 8'hFC;
			14'd10712: ff_rdata <= 8'h69;
			14'd10713: ff_rdata <= 8'hE1;
			14'd10714: ff_rdata <= 8'hC9;
			14'd10715: ff_rdata <= 8'h79;
			14'd10716: ff_rdata <= 8'hE6;
			14'd10717: ff_rdata <= 8'h1F;
			14'd10718: ff_rdata <= 8'hC8;
			14'd10719: ff_rdata <= 8'hE5;
			14'd10720: ff_rdata <= 8'hC5;
			14'd10721: ff_rdata <= 8'h21;
			14'd10722: ff_rdata <= 8'hB7;
			14'd10723: ff_rdata <= 8'hFA;
			14'd10724: ff_rdata <= 8'h57;
			14'd10725: ff_rdata <= 8'h7B;
			14'd10726: ff_rdata <= 8'h0F;
			14'd10727: ff_rdata <= 8'h0F;
			14'd10728: ff_rdata <= 8'h0F;
			14'd10729: ff_rdata <= 8'hE6;
			14'd10730: ff_rdata <= 8'h07;
			14'd10731: ff_rdata <= 8'h5F;
			14'd10732: ff_rdata <= 8'h06;
			14'd10733: ff_rdata <= 8'h05;
			14'd10734: ff_rdata <= 8'hCB;
			14'd10735: ff_rdata <= 8'h1A;
			14'd10736: ff_rdata <= 8'h30;
			14'd10737: ff_rdata <= 8'h01;
			14'd10738: ff_rdata <= 8'h73;
			14'd10739: ff_rdata <= 8'h23;
			14'd10740: ff_rdata <= 8'h10;
			14'd10741: ff_rdata <= 8'hF8;
			14'd10742: ff_rdata <= 8'hCD;
			14'd10743: ff_rdata <= 8'hFC;
			14'd10744: ff_rdata <= 8'h69;
			14'd10745: ff_rdata <= 8'hC1;
			14'd10746: ff_rdata <= 8'hE1;
			14'd10747: ff_rdata <= 8'hC9;
			14'd10748: ff_rdata <= 8'h21;
			14'd10749: ff_rdata <= 8'hB7;
			14'd10750: ff_rdata <= 8'hFA;
			14'd10751: ff_rdata <= 8'h3A;
			14'd10752: ff_rdata <= 8'h89;
			14'd10753: ff_rdata <= 8'hFA;
			14'd10754: ff_rdata <= 8'h57;
			14'd10755: ff_rdata <= 8'h86;
			14'd10756: ff_rdata <= 8'h23;
			14'd10757: ff_rdata <= 8'h07;
			14'd10758: ff_rdata <= 8'h07;
			14'd10759: ff_rdata <= 8'h07;
			14'd10760: ff_rdata <= 8'h07;
			14'd10761: ff_rdata <= 8'h47;
			14'd10762: ff_rdata <= 8'h0E;
			14'd10763: ff_rdata <= 8'h37;
			14'd10764: ff_rdata <= 8'hCD;
			14'd10765: ff_rdata <= 8'h36;
			14'd10766: ff_rdata <= 8'h6A;
			14'd10767: ff_rdata <= 8'h7A;
			14'd10768: ff_rdata <= 8'h86;
			14'd10769: ff_rdata <= 8'h23;
			14'd10770: ff_rdata <= 8'h47;
			14'd10771: ff_rdata <= 8'h0E;
			14'd10772: ff_rdata <= 8'h38;
			14'd10773: ff_rdata <= 8'hCD;
			14'd10774: ff_rdata <= 8'h40;
			14'd10775: ff_rdata <= 8'h6A;
			14'd10776: ff_rdata <= 8'h7A;
			14'd10777: ff_rdata <= 8'h86;
			14'd10778: ff_rdata <= 8'h23;
			14'd10779: ff_rdata <= 8'h07;
			14'd10780: ff_rdata <= 8'h07;
			14'd10781: ff_rdata <= 8'h07;
			14'd10782: ff_rdata <= 8'h07;
			14'd10783: ff_rdata <= 8'h47;
			14'd10784: ff_rdata <= 8'hCD;
			14'd10785: ff_rdata <= 8'h36;
			14'd10786: ff_rdata <= 8'h6A;
			14'd10787: ff_rdata <= 8'h7A;
			14'd10788: ff_rdata <= 8'h86;
			14'd10789: ff_rdata <= 8'h23;
			14'd10790: ff_rdata <= 8'h47;
			14'd10791: ff_rdata <= 8'h0E;
			14'd10792: ff_rdata <= 8'h37;
			14'd10793: ff_rdata <= 8'hCD;
			14'd10794: ff_rdata <= 8'h40;
			14'd10795: ff_rdata <= 8'h6A;
			14'd10796: ff_rdata <= 8'h7A;
			14'd10797: ff_rdata <= 8'h86;
			14'd10798: ff_rdata <= 8'h23;
			14'd10799: ff_rdata <= 8'h47;
			14'd10800: ff_rdata <= 8'h0E;
			14'd10801: ff_rdata <= 8'h36;
			14'd10802: ff_rdata <= 8'hCD;
			14'd10803: ff_rdata <= 8'h40;
			14'd10804: ff_rdata <= 8'h6A;
			14'd10805: ff_rdata <= 8'hC9;
			14'd10806: ff_rdata <= 8'hCD;
			14'd10807: ff_rdata <= 8'hE0;
			14'd10808: ff_rdata <= 8'h6D;
			14'd10809: ff_rdata <= 8'hE6;
			14'd10810: ff_rdata <= 8'h0F;
			14'd10811: ff_rdata <= 8'hB0;
			14'd10812: ff_rdata <= 8'h47;
			14'd10813: ff_rdata <= 8'hC3;
			14'd10814: ff_rdata <= 8'hB5;
			14'd10815: ff_rdata <= 8'h6D;
			14'd10816: ff_rdata <= 8'hCD;
			14'd10817: ff_rdata <= 8'hE0;
			14'd10818: ff_rdata <= 8'h6D;
			14'd10819: ff_rdata <= 8'hE6;
			14'd10820: ff_rdata <= 8'hF0;
			14'd10821: ff_rdata <= 8'h18;
			14'd10822: ff_rdata <= 8'hF4;
			14'd10823: ff_rdata <= 8'hC3;
			14'd10824: ff_rdata <= 8'h58;
			14'd10825: ff_rdata <= 8'h6C;
			14'd10826: ff_rdata <= 8'hC5;
			14'd10827: ff_rdata <= 8'hD5;
			14'd10828: ff_rdata <= 8'hCD;
			14'd10829: ff_rdata <= 8'h58;
			14'd10830: ff_rdata <= 8'h6C;
			14'd10831: ff_rdata <= 8'hD1;
			14'd10832: ff_rdata <= 8'hC1;
			14'd10833: ff_rdata <= 8'h3E;
			14'd10834: ff_rdata <= 8'h0F;
			14'd10835: ff_rdata <= 8'h91;
			14'd10836: ff_rdata <= 8'h0F;
			14'd10837: ff_rdata <= 8'hE6;
			14'd10838: ff_rdata <= 8'h07;
			14'd10839: ff_rdata <= 8'hDD;
			14'd10840: ff_rdata <= 8'h77;
			14'd10841: ff_rdata <= 8'h01;
			14'd10842: ff_rdata <= 8'hCB;
			14'd10843: ff_rdata <= 8'hBA;
			14'd10844: ff_rdata <= 8'hDD;
			14'd10845: ff_rdata <= 8'h73;
			14'd10846: ff_rdata <= 8'h03;
			14'd10847: ff_rdata <= 8'hDD;
			14'd10848: ff_rdata <= 8'h72;
			14'd10849: ff_rdata <= 8'h04;
			14'd10850: ff_rdata <= 8'hCD;
			14'd10851: ff_rdata <= 8'h78;
			14'd10852: ff_rdata <= 8'h6A;
			14'd10853: ff_rdata <= 8'hCD;
			14'd10854: ff_rdata <= 8'h3A;
			14'd10855: ff_rdata <= 8'h6C;
			14'd10856: ff_rdata <= 8'hDD;
			14'd10857: ff_rdata <= 8'h7E;
			14'd10858: ff_rdata <= 8'h00;
			14'd10859: ff_rdata <= 8'hC6;
			14'd10860: ff_rdata <= 8'h10;
			14'd10861: ff_rdata <= 8'h4F;
			14'd10862: ff_rdata <= 8'hCD;
			14'd10863: ff_rdata <= 8'hE0;
			14'd10864: ff_rdata <= 8'h6D;
			14'd10865: ff_rdata <= 8'hF6;
			14'd10866: ff_rdata <= 8'h10;
			14'd10867: ff_rdata <= 8'h47;
			14'd10868: ff_rdata <= 8'hCD;
			14'd10869: ff_rdata <= 8'hB5;
			14'd10870: ff_rdata <= 8'h6D;
			14'd10871: ff_rdata <= 8'hC9;
			14'd10872: ff_rdata <= 8'hDD;
			14'd10873: ff_rdata <= 8'h6E;
			14'd10874: ff_rdata <= 8'h05;
			14'd10875: ff_rdata <= 8'hDD;
			14'd10876: ff_rdata <= 8'h66;
			14'd10877: ff_rdata <= 8'h06;
			14'd10878: ff_rdata <= 8'hDD;
			14'd10879: ff_rdata <= 8'h5E;
			14'd10880: ff_rdata <= 8'h03;
			14'd10881: ff_rdata <= 8'hDD;
			14'd10882: ff_rdata <= 8'h56;
			14'd10883: ff_rdata <= 8'h04;
			14'd10884: ff_rdata <= 8'h19;
			14'd10885: ff_rdata <= 8'hDD;
			14'd10886: ff_rdata <= 8'h5E;
			14'd10887: ff_rdata <= 8'h07;
			14'd10888: ff_rdata <= 8'hDD;
			14'd10889: ff_rdata <= 8'h56;
			14'd10890: ff_rdata <= 8'h08;
			14'd10891: ff_rdata <= 8'h19;
			14'd10892: ff_rdata <= 8'h11;
			14'd10893: ff_rdata <= 8'h29;
			14'd10894: ff_rdata <= 8'h05;
			14'd10895: ff_rdata <= 8'h19;
			14'd10896: ff_rdata <= 8'h7C;
			14'd10897: ff_rdata <= 8'hA7;
			14'd10898: ff_rdata <= 8'hF2;
			14'd10899: ff_rdata <= 8'hA5;
			14'd10900: ff_rdata <= 8'h6A;
			14'd10901: ff_rdata <= 8'hFE;
			14'd10902: ff_rdata <= 8'hC4;
			14'd10903: ff_rdata <= 8'h30;
			14'd10904: ff_rdata <= 8'h07;
			14'd10905: ff_rdata <= 8'hD6;
			14'd10906: ff_rdata <= 8'h0C;
			14'd10907: ff_rdata <= 8'hFA;
			14'd10908: ff_rdata <= 8'h99;
			14'd10909: ff_rdata <= 8'h6A;
			14'd10910: ff_rdata <= 8'h18;
			14'd10911: ff_rdata <= 8'h05;
			14'd10912: ff_rdata <= 8'hC6;
			14'd10913: ff_rdata <= 8'h0C;
			14'd10914: ff_rdata <= 8'hFA;
			14'd10915: ff_rdata <= 8'hA0;
			14'd10916: ff_rdata <= 8'h6A;
			14'd10917: ff_rdata <= 8'h67;
			14'd10918: ff_rdata <= 8'h4D;
			14'd10919: ff_rdata <= 8'h2E;
			14'd10920: ff_rdata <= 8'h00;
			14'd10921: ff_rdata <= 8'h11;
			14'd10922: ff_rdata <= 8'h04;
			14'd10923: ff_rdata <= 8'hF4;
			14'd10924: ff_rdata <= 8'hD6;
			14'd10925: ff_rdata <= 8'h3C;
			14'd10926: ff_rdata <= 8'h38;
			14'd10927: ff_rdata <= 8'h03;
			14'd10928: ff_rdata <= 8'h67;
			14'd10929: ff_rdata <= 8'h2E;
			14'd10930: ff_rdata <= 8'h14;
			14'd10931: ff_rdata <= 8'h19;
			14'd10932: ff_rdata <= 8'hDA;
			14'd10933: ff_rdata <= 8'hB3;
			14'd10934: ff_rdata <= 8'h6A;
			14'd10935: ff_rdata <= 8'hED;
			14'd10936: ff_rdata <= 8'h52;
			14'd10937: ff_rdata <= 8'h45;
			14'd10938: ff_rdata <= 8'h7C;
			14'd10939: ff_rdata <= 8'h84;
			14'd10940: ff_rdata <= 8'h84;
			14'd10941: ff_rdata <= 8'h21;
			14'd10942: ff_rdata <= 8'h2C;
			14'd10943: ff_rdata <= 8'h6B;
			14'd10944: ff_rdata <= 8'hCD;
			14'd10945: ff_rdata <= 8'h86;
			14'd10946: ff_rdata <= 8'h54;
			14'd10947: ff_rdata <= 8'h78;
			14'd10948: ff_rdata <= 8'h5E;
			14'd10949: ff_rdata <= 8'h23;
			14'd10950: ff_rdata <= 8'h56;
			14'd10951: ff_rdata <= 8'h23;
			14'd10952: ff_rdata <= 8'h66;
			14'd10953: ff_rdata <= 8'h2E;
			14'd10954: ff_rdata <= 8'h00;
			14'd10955: ff_rdata <= 8'h45;
			14'd10956: ff_rdata <= 8'h29;
			14'd10957: ff_rdata <= 8'h30;
			14'd10958: ff_rdata <= 8'h01;
			14'd10959: ff_rdata <= 8'h09;
			14'd10960: ff_rdata <= 8'h29;
			14'd10961: ff_rdata <= 8'h30;
			14'd10962: ff_rdata <= 8'h01;
			14'd10963: ff_rdata <= 8'h09;
			14'd10964: ff_rdata <= 8'h29;
			14'd10965: ff_rdata <= 8'h30;
			14'd10966: ff_rdata <= 8'h01;
			14'd10967: ff_rdata <= 8'h09;
			14'd10968: ff_rdata <= 8'h29;
			14'd10969: ff_rdata <= 8'h30;
			14'd10970: ff_rdata <= 8'h01;
			14'd10971: ff_rdata <= 8'h09;
			14'd10972: ff_rdata <= 8'h29;
			14'd10973: ff_rdata <= 8'h30;
			14'd10974: ff_rdata <= 8'h01;
			14'd10975: ff_rdata <= 8'h09;
			14'd10976: ff_rdata <= 8'h29;
			14'd10977: ff_rdata <= 8'h30;
			14'd10978: ff_rdata <= 8'h01;
			14'd10979: ff_rdata <= 8'h09;
			14'd10980: ff_rdata <= 8'h29;
			14'd10981: ff_rdata <= 8'h30;
			14'd10982: ff_rdata <= 8'h01;
			14'd10983: ff_rdata <= 8'h09;
			14'd10984: ff_rdata <= 8'h29;
			14'd10985: ff_rdata <= 8'h30;
			14'd10986: ff_rdata <= 8'h01;
			14'd10987: ff_rdata <= 8'h09;
			14'd10988: ff_rdata <= 8'h6C;
			14'd10989: ff_rdata <= 8'h60;
			14'd10990: ff_rdata <= 8'h19;
			14'd10991: ff_rdata <= 8'hCB;
			14'd10992: ff_rdata <= 8'h3C;
			14'd10993: ff_rdata <= 8'hCB;
			14'd10994: ff_rdata <= 8'h1D;
			14'd10995: ff_rdata <= 8'hCB;
			14'd10996: ff_rdata <= 8'h3C;
			14'd10997: ff_rdata <= 8'hCB;
			14'd10998: ff_rdata <= 8'h1D;
			14'd10999: ff_rdata <= 8'h30;
			14'd11000: ff_rdata <= 8'h06;
			14'd11001: ff_rdata <= 8'h23;
			14'd11002: ff_rdata <= 8'hCB;
			14'd11003: ff_rdata <= 8'h54;
			14'd11004: ff_rdata <= 8'h28;
			14'd11005: ff_rdata <= 8'h01;
			14'd11006: ff_rdata <= 8'h2B;
			14'd11007: ff_rdata <= 8'hD6;
			14'd11008: ff_rdata <= 8'h08;
			14'd11009: ff_rdata <= 8'h30;
			14'd11010: ff_rdata <= 8'h08;
			14'd11011: ff_rdata <= 8'hCB;
			14'd11012: ff_rdata <= 8'h3C;
			14'd11013: ff_rdata <= 8'hCB;
			14'd11014: ff_rdata <= 8'h1D;
			14'd11015: ff_rdata <= 8'hC6;
			14'd11016: ff_rdata <= 8'h04;
			14'd11017: ff_rdata <= 8'h20;
			14'd11018: ff_rdata <= 8'hF8;
			14'd11019: ff_rdata <= 8'hFE;
			14'd11020: ff_rdata <= 8'h20;
			14'd11021: ff_rdata <= 8'h38;
			14'd11022: ff_rdata <= 8'h02;
			14'd11023: ff_rdata <= 8'h3E;
			14'd11024: ff_rdata <= 8'h1C;
			14'd11025: ff_rdata <= 8'hB4;
			14'd11026: ff_rdata <= 8'h1F;
			14'd11027: ff_rdata <= 8'h67;
			14'd11028: ff_rdata <= 8'hCB;
			14'd11029: ff_rdata <= 8'h1D;
			14'd11030: ff_rdata <= 8'hDD;
			14'd11031: ff_rdata <= 8'h4E;
			14'd11032: ff_rdata <= 8'h00;
			14'd11033: ff_rdata <= 8'h45;
			14'd11034: ff_rdata <= 8'hCD;
			14'd11035: ff_rdata <= 8'hB5;
			14'd11036: ff_rdata <= 8'h6D;
			14'd11037: ff_rdata <= 8'h79;
			14'd11038: ff_rdata <= 8'hC6;
			14'd11039: ff_rdata <= 8'h10;
			14'd11040: ff_rdata <= 8'h4F;
			14'd11041: ff_rdata <= 8'hCD;
			14'd11042: ff_rdata <= 8'hE0;
			14'd11043: ff_rdata <= 8'h6D;
			14'd11044: ff_rdata <= 8'hE6;
			14'd11045: ff_rdata <= 8'h30;
			14'd11046: ff_rdata <= 8'hB4;
			14'd11047: ff_rdata <= 8'h47;
			14'd11048: ff_rdata <= 8'hCD;
			14'd11049: ff_rdata <= 8'hB5;
			14'd11050: ff_rdata <= 8'h6D;
			14'd11051: ff_rdata <= 8'hC9;
			14'd11052: ff_rdata <= 8'h00;
			14'd11053: ff_rdata <= 8'h08;
			14'd11054: ff_rdata <= 8'h79;
			14'd11055: ff_rdata <= 8'h79;
			14'd11056: ff_rdata <= 8'h08;
			14'd11057: ff_rdata <= 8'h81;
			14'd11058: ff_rdata <= 8'hFA;
			14'd11059: ff_rdata <= 8'h08;
			14'd11060: ff_rdata <= 8'h89;
			14'd11061: ff_rdata <= 8'h83;
			14'd11062: ff_rdata <= 8'h09;
			14'd11063: ff_rdata <= 8'h91;
			14'd11064: ff_rdata <= 8'h14;
			14'd11065: ff_rdata <= 8'h0A;
			14'd11066: ff_rdata <= 8'h99;
			14'd11067: ff_rdata <= 8'hAD;
			14'd11068: ff_rdata <= 8'h0A;
			14'd11069: ff_rdata <= 8'hA3;
			14'd11070: ff_rdata <= 8'h50;
			14'd11071: ff_rdata <= 8'h0B;
			14'd11072: ff_rdata <= 8'hAC;
			14'd11073: ff_rdata <= 8'hFC;
			14'd11074: ff_rdata <= 8'h0B;
			14'd11075: ff_rdata <= 8'hB6;
			14'd11076: ff_rdata <= 8'hB2;
			14'd11077: ff_rdata <= 8'h0C;
			14'd11078: ff_rdata <= 8'hC2;
			14'd11079: ff_rdata <= 8'h74;
			14'd11080: ff_rdata <= 8'h0D;
			14'd11081: ff_rdata <= 8'hCD;
			14'd11082: ff_rdata <= 8'h41;
			14'd11083: ff_rdata <= 8'h0E;
			14'd11084: ff_rdata <= 8'hD9;
			14'd11085: ff_rdata <= 8'h1A;
			14'd11086: ff_rdata <= 8'h0F;
			14'd11087: ff_rdata <= 8'hE6;
			14'd11088: ff_rdata <= 8'h50;
			14'd11089: ff_rdata <= 8'h59;
			14'd11090: ff_rdata <= 8'hCD;
			14'd11091: ff_rdata <= 8'h62;
			14'd11092: ff_rdata <= 8'h6B;
			14'd11093: ff_rdata <= 8'hD8;
			14'd11094: ff_rdata <= 8'hED;
			14'd11095: ff_rdata <= 8'h53;
			14'd11096: ff_rdata <= 8'h9D;
			14'd11097: ff_rdata <= 8'hF9;
			14'd11098: ff_rdata <= 8'h2A;
			14'd11099: ff_rdata <= 8'h9F;
			14'd11100: ff_rdata <= 8'hF9;
			14'd11101: ff_rdata <= 8'h19;
			14'd11102: ff_rdata <= 8'hEB;
			14'd11103: ff_rdata <= 8'hC3;
			14'd11104: ff_rdata <= 8'hE9;
			14'd11105: ff_rdata <= 8'h6B;
			14'd11106: ff_rdata <= 8'h21;
			14'd11107: ff_rdata <= 8'h34;
			14'd11108: ff_rdata <= 8'hFE;
			14'd11109: ff_rdata <= 8'h19;
			14'd11110: ff_rdata <= 8'hD8;
			14'd11111: ff_rdata <= 8'h21;
			14'd11112: ff_rdata <= 8'h66;
			14'd11113: ff_rdata <= 8'hFE;
			14'd11114: ff_rdata <= 8'h19;
			14'd11115: ff_rdata <= 8'h3F;
			14'd11116: ff_rdata <= 8'hD8;
			14'd11117: ff_rdata <= 8'h29;
			14'd11118: ff_rdata <= 8'h11;
			14'd11119: ff_rdata <= 8'h76;
			14'd11120: ff_rdata <= 8'h6B;
			14'd11121: ff_rdata <= 8'h19;
			14'd11122: ff_rdata <= 8'h5E;
			14'd11123: ff_rdata <= 8'h23;
			14'd11124: ff_rdata <= 8'h56;
			14'd11125: ff_rdata <= 8'hC9;
			14'd11126: ff_rdata <= 8'hC7;
			14'd11127: ff_rdata <= 8'hFE;
			14'd11128: ff_rdata <= 8'hD2;
			14'd11129: ff_rdata <= 8'hFE;
			14'd11130: ff_rdata <= 8'hDD;
			14'd11131: ff_rdata <= 8'hFE;
			14'd11132: ff_rdata <= 8'hE7;
			14'd11133: ff_rdata <= 8'hFE;
			14'd11134: ff_rdata <= 8'hF2;
			14'd11135: ff_rdata <= 8'hFE;
			14'd11136: ff_rdata <= 8'hFD;
			14'd11137: ff_rdata <= 8'hFE;
			14'd11138: ff_rdata <= 8'h07;
			14'd11139: ff_rdata <= 8'hFF;
			14'd11140: ff_rdata <= 8'h12;
			14'd11141: ff_rdata <= 8'hFF;
			14'd11142: ff_rdata <= 8'h1D;
			14'd11143: ff_rdata <= 8'hFF;
			14'd11144: ff_rdata <= 8'h27;
			14'd11145: ff_rdata <= 8'hFF;
			14'd11146: ff_rdata <= 8'h32;
			14'd11147: ff_rdata <= 8'hFF;
			14'd11148: ff_rdata <= 8'h3C;
			14'd11149: ff_rdata <= 8'hFF;
			14'd11150: ff_rdata <= 8'h47;
			14'd11151: ff_rdata <= 8'hFF;
			14'd11152: ff_rdata <= 8'h51;
			14'd11153: ff_rdata <= 8'hFF;
			14'd11154: ff_rdata <= 8'h5C;
			14'd11155: ff_rdata <= 8'hFF;
			14'd11156: ff_rdata <= 8'h66;
			14'd11157: ff_rdata <= 8'hFF;
			14'd11158: ff_rdata <= 8'h71;
			14'd11159: ff_rdata <= 8'hFF;
			14'd11160: ff_rdata <= 8'h7B;
			14'd11161: ff_rdata <= 8'hFF;
			14'd11162: ff_rdata <= 8'h85;
			14'd11163: ff_rdata <= 8'hFF;
			14'd11164: ff_rdata <= 8'h90;
			14'd11165: ff_rdata <= 8'hFF;
			14'd11166: ff_rdata <= 8'h9A;
			14'd11167: ff_rdata <= 8'hFF;
			14'd11168: ff_rdata <= 8'hA4;
			14'd11169: ff_rdata <= 8'hFF;
			14'd11170: ff_rdata <= 8'hAF;
			14'd11171: ff_rdata <= 8'hFF;
			14'd11172: ff_rdata <= 8'hB9;
			14'd11173: ff_rdata <= 8'hFF;
			14'd11174: ff_rdata <= 8'hC3;
			14'd11175: ff_rdata <= 8'hFF;
			14'd11176: ff_rdata <= 8'hCD;
			14'd11177: ff_rdata <= 8'hFF;
			14'd11178: ff_rdata <= 8'hD8;
			14'd11179: ff_rdata <= 8'hFF;
			14'd11180: ff_rdata <= 8'hE2;
			14'd11181: ff_rdata <= 8'hFF;
			14'd11182: ff_rdata <= 8'hEC;
			14'd11183: ff_rdata <= 8'hFF;
			14'd11184: ff_rdata <= 8'hF6;
			14'd11185: ff_rdata <= 8'hFF;
			14'd11186: ff_rdata <= 8'h00;
			14'd11187: ff_rdata <= 8'h00;
			14'd11188: ff_rdata <= 8'h0A;
			14'd11189: ff_rdata <= 8'h00;
			14'd11190: ff_rdata <= 8'h14;
			14'd11191: ff_rdata <= 8'h00;
			14'd11192: ff_rdata <= 8'h1E;
			14'd11193: ff_rdata <= 8'h00;
			14'd11194: ff_rdata <= 8'h28;
			14'd11195: ff_rdata <= 8'h00;
			14'd11196: ff_rdata <= 8'h32;
			14'd11197: ff_rdata <= 8'h00;
			14'd11198: ff_rdata <= 8'h3C;
			14'd11199: ff_rdata <= 8'h00;
			14'd11200: ff_rdata <= 8'h46;
			14'd11201: ff_rdata <= 8'h00;
			14'd11202: ff_rdata <= 8'h50;
			14'd11203: ff_rdata <= 8'h00;
			14'd11204: ff_rdata <= 8'h5A;
			14'd11205: ff_rdata <= 8'h00;
			14'd11206: ff_rdata <= 8'h64;
			14'd11207: ff_rdata <= 8'h00;
			14'd11208: ff_rdata <= 8'h6D;
			14'd11209: ff_rdata <= 8'h00;
			14'd11210: ff_rdata <= 8'h77;
			14'd11211: ff_rdata <= 8'h00;
			14'd11212: ff_rdata <= 8'h81;
			14'd11213: ff_rdata <= 8'h00;
			14'd11214: ff_rdata <= 8'h8B;
			14'd11215: ff_rdata <= 8'h00;
			14'd11216: ff_rdata <= 8'h95;
			14'd11217: ff_rdata <= 8'h00;
			14'd11218: ff_rdata <= 8'h9E;
			14'd11219: ff_rdata <= 8'h00;
			14'd11220: ff_rdata <= 8'hA8;
			14'd11221: ff_rdata <= 8'h00;
			14'd11222: ff_rdata <= 8'hB2;
			14'd11223: ff_rdata <= 8'h00;
			14'd11224: ff_rdata <= 8'hBB;
			14'd11225: ff_rdata <= 8'h00;
			14'd11226: ff_rdata <= 8'h50;
			14'd11227: ff_rdata <= 8'h59;
			14'd11228: ff_rdata <= 8'hCD;
			14'd11229: ff_rdata <= 8'h0F;
			14'd11230: ff_rdata <= 8'h6C;
			14'd11231: ff_rdata <= 8'hD8;
			14'd11232: ff_rdata <= 8'hED;
			14'd11233: ff_rdata <= 8'h53;
			14'd11234: ff_rdata <= 8'h9F;
			14'd11235: ff_rdata <= 8'hF9;
			14'd11236: ff_rdata <= 8'h2A;
			14'd11237: ff_rdata <= 8'h9D;
			14'd11238: ff_rdata <= 8'hF9;
			14'd11239: ff_rdata <= 8'h19;
			14'd11240: ff_rdata <= 8'hEB;
			14'd11241: ff_rdata <= 8'hDD;
			14'd11242: ff_rdata <= 8'h21;
			14'd11243: ff_rdata <= 8'h27;
			14'd11244: ff_rdata <= 8'hFA;
			14'd11245: ff_rdata <= 8'h06;
			14'd11246: ff_rdata <= 8'h09;
			14'd11247: ff_rdata <= 8'h0E;
			14'd11248: ff_rdata <= 8'h0E;
			14'd11249: ff_rdata <= 8'hCD;
			14'd11250: ff_rdata <= 8'hE0;
			14'd11251: ff_rdata <= 8'h6D;
			14'd11252: ff_rdata <= 8'hE6;
			14'd11253: ff_rdata <= 8'h20;
			14'd11254: ff_rdata <= 8'h28;
			14'd11255: ff_rdata <= 8'h02;
			14'd11256: ff_rdata <= 8'h06;
			14'd11257: ff_rdata <= 8'h06;
			14'd11258: ff_rdata <= 8'hC5;
			14'd11259: ff_rdata <= 8'hD5;
			14'd11260: ff_rdata <= 8'hDD;
			14'd11261: ff_rdata <= 8'h73;
			14'd11262: ff_rdata <= 8'h05;
			14'd11263: ff_rdata <= 8'hDD;
			14'd11264: ff_rdata <= 8'h72;
			14'd11265: ff_rdata <= 8'h06;
			14'd11266: ff_rdata <= 8'hCD;
			14'd11267: ff_rdata <= 8'h78;
			14'd11268: ff_rdata <= 8'h6A;
			14'd11269: ff_rdata <= 8'h01;
			14'd11270: ff_rdata <= 8'h10;
			14'd11271: ff_rdata <= 8'h00;
			14'd11272: ff_rdata <= 8'hDD;
			14'd11273: ff_rdata <= 8'h09;
			14'd11274: ff_rdata <= 8'hD1;
			14'd11275: ff_rdata <= 8'hC1;
			14'd11276: ff_rdata <= 8'h10;
			14'd11277: ff_rdata <= 8'hEC;
			14'd11278: ff_rdata <= 8'hC9;
			14'd11279: ff_rdata <= 8'h7A;
			14'd11280: ff_rdata <= 8'hA7;
			14'd11281: ff_rdata <= 8'hF5;
			14'd11282: ff_rdata <= 8'hFC;
			14'd11283: ff_rdata <= 8'h32;
			14'd11284: ff_rdata <= 8'h6C;
			14'd11285: ff_rdata <= 8'h7A;
			14'd11286: ff_rdata <= 8'h63;
			14'd11287: ff_rdata <= 8'h2E;
			14'd11288: ff_rdata <= 8'h00;
			14'd11289: ff_rdata <= 8'h11;
			14'd11290: ff_rdata <= 8'h0F;
			14'd11291: ff_rdata <= 8'h64;
			14'd11292: ff_rdata <= 8'h29;
			14'd11293: ff_rdata <= 8'h17;
			14'd11294: ff_rdata <= 8'hBA;
			14'd11295: ff_rdata <= 8'h38;
			14'd11296: ff_rdata <= 8'h03;
			14'd11297: ff_rdata <= 8'hF1;
			14'd11298: ff_rdata <= 8'h37;
			14'd11299: ff_rdata <= 8'hC9;
			14'd11300: ff_rdata <= 8'h29;
			14'd11301: ff_rdata <= 8'h17;
			14'd11302: ff_rdata <= 8'hBA;
			14'd11303: ff_rdata <= 8'h38;
			14'd11304: ff_rdata <= 8'h02;
			14'd11305: ff_rdata <= 8'h92;
			14'd11306: ff_rdata <= 8'h2C;
			14'd11307: ff_rdata <= 8'h1D;
			14'd11308: ff_rdata <= 8'hC2;
			14'd11309: ff_rdata <= 8'h24;
			14'd11310: ff_rdata <= 8'h6C;
			14'd11311: ff_rdata <= 8'hEB;
			14'd11312: ff_rdata <= 8'hF1;
			14'd11313: ff_rdata <= 8'hF0;
			14'd11314: ff_rdata <= 8'hAF;
			14'd11315: ff_rdata <= 8'h67;
			14'd11316: ff_rdata <= 8'h6F;
			14'd11317: ff_rdata <= 8'hED;
			14'd11318: ff_rdata <= 8'h52;
			14'd11319: ff_rdata <= 8'hEB;
			14'd11320: ff_rdata <= 8'hA7;
			14'd11321: ff_rdata <= 8'hC9;
			14'd11322: ff_rdata <= 8'hDD;
			14'd11323: ff_rdata <= 8'h7E;
			14'd11324: ff_rdata <= 8'h02;
			14'd11325: ff_rdata <= 8'hDD;
			14'd11326: ff_rdata <= 8'h86;
			14'd11327: ff_rdata <= 8'h01;
			14'd11328: ff_rdata <= 8'hFE;
			14'd11329: ff_rdata <= 8'h10;
			14'd11330: ff_rdata <= 8'h38;
			14'd11331: ff_rdata <= 8'h02;
			14'd11332: ff_rdata <= 8'h3E;
			14'd11333: ff_rdata <= 8'h0F;
			14'd11334: ff_rdata <= 8'h47;
			14'd11335: ff_rdata <= 8'hDD;
			14'd11336: ff_rdata <= 8'h7E;
			14'd11337: ff_rdata <= 8'h00;
			14'd11338: ff_rdata <= 8'hC6;
			14'd11339: ff_rdata <= 8'h20;
			14'd11340: ff_rdata <= 8'h4F;
			14'd11341: ff_rdata <= 8'hCD;
			14'd11342: ff_rdata <= 8'hE0;
			14'd11343: ff_rdata <= 8'h6D;
			14'd11344: ff_rdata <= 8'hE6;
			14'd11345: ff_rdata <= 8'hF0;
			14'd11346: ff_rdata <= 8'hB0;
			14'd11347: ff_rdata <= 8'h47;
			14'd11348: ff_rdata <= 8'hCD;
			14'd11349: ff_rdata <= 8'hB5;
			14'd11350: ff_rdata <= 8'h6D;
			14'd11351: ff_rdata <= 8'hC9;
			14'd11352: ff_rdata <= 8'hDD;
			14'd11353: ff_rdata <= 8'h7E;
			14'd11354: ff_rdata <= 8'h00;
			14'd11355: ff_rdata <= 8'hC6;
			14'd11356: ff_rdata <= 8'h10;
			14'd11357: ff_rdata <= 8'h4F;
			14'd11358: ff_rdata <= 8'hCD;
			14'd11359: ff_rdata <= 8'hE0;
			14'd11360: ff_rdata <= 8'h6D;
			14'd11361: ff_rdata <= 8'hE6;
			14'd11362: ff_rdata <= 8'h2F;
			14'd11363: ff_rdata <= 8'h47;
			14'd11364: ff_rdata <= 8'hCD;
			14'd11365: ff_rdata <= 8'hB5;
			14'd11366: ff_rdata <= 8'h6D;
			14'd11367: ff_rdata <= 8'hC9;
			14'd11368: ff_rdata <= 8'hE5;
			14'd11369: ff_rdata <= 8'h79;
			14'd11370: ff_rdata <= 8'hE6;
			14'd11371: ff_rdata <= 8'h1F;
			14'd11372: ff_rdata <= 8'h57;
			14'd11373: ff_rdata <= 8'h2F;
			14'd11374: ff_rdata <= 8'h5F;
			14'd11375: ff_rdata <= 8'h0E;
			14'd11376: ff_rdata <= 8'h0E;
			14'd11377: ff_rdata <= 8'hCD;
			14'd11378: ff_rdata <= 8'hE0;
			14'd11379: ff_rdata <= 8'h6D;
			14'd11380: ff_rdata <= 8'h6F;
			14'd11381: ff_rdata <= 8'hA3;
			14'd11382: ff_rdata <= 8'h47;
			14'd11383: ff_rdata <= 8'hCD;
			14'd11384: ff_rdata <= 8'hB5;
			14'd11385: ff_rdata <= 8'h6D;
			14'd11386: ff_rdata <= 8'h7D;
			14'd11387: ff_rdata <= 8'hB2;
			14'd11388: ff_rdata <= 8'h47;
			14'd11389: ff_rdata <= 8'hCD;
			14'd11390: ff_rdata <= 8'hB5;
			14'd11391: ff_rdata <= 8'h6D;
			14'd11392: ff_rdata <= 8'hE1;
			14'd11393: ff_rdata <= 8'hC9;
			14'd11394: ff_rdata <= 8'hE5;
			14'd11395: ff_rdata <= 8'h7A;
			14'd11396: ff_rdata <= 8'hD6;
			14'd11397: ff_rdata <= 8'h3C;
			14'd11398: ff_rdata <= 8'h26;
			14'd11399: ff_rdata <= 8'h0C;
			14'd11400: ff_rdata <= 8'h38;
			14'd11401: ff_rdata <= 8'h04;
			14'd11402: ff_rdata <= 8'h94;
			14'd11403: ff_rdata <= 8'hD2;
			14'd11404: ff_rdata <= 8'h8A;
			14'd11405: ff_rdata <= 8'h6C;
			14'd11406: ff_rdata <= 8'h84;
			14'd11407: ff_rdata <= 8'hD2;
			14'd11408: ff_rdata <= 8'h8E;
			14'd11409: ff_rdata <= 8'h6C;
			14'd11410: ff_rdata <= 8'h2A;
			14'd11411: ff_rdata <= 8'hA1;
			14'd11412: ff_rdata <= 8'hF9;
			14'd11413: ff_rdata <= 8'hCD;
			14'd11414: ff_rdata <= 8'h86;
			14'd11415: ff_rdata <= 8'h54;
			14'd11416: ff_rdata <= 8'h5E;
			14'd11417: ff_rdata <= 8'hE1;
			14'd11418: ff_rdata <= 8'hCB;
			14'd11419: ff_rdata <= 8'h7B;
			14'd11420: ff_rdata <= 8'hC8;
			14'd11421: ff_rdata <= 8'h15;
			14'd11422: ff_rdata <= 8'hC9;
			14'd11423: ff_rdata <= 8'h79;
			14'd11424: ff_rdata <= 8'hFE;
			14'd11425: ff_rdata <= 8'h16;
			14'd11426: ff_rdata <= 8'h3F;
			14'd11427: ff_rdata <= 8'hD8;
			14'd11428: ff_rdata <= 8'hE5;
			14'd11429: ff_rdata <= 8'hFE;
			14'd11430: ff_rdata <= 8'h0A;
			14'd11431: ff_rdata <= 8'h38;
			14'd11432: ff_rdata <= 8'h04;
			14'd11433: ff_rdata <= 8'hC6;
			14'd11434: ff_rdata <= 8'h6E;
			14'd11435: ff_rdata <= 8'h18;
			14'd11436: ff_rdata <= 8'h05;
			14'd11437: ff_rdata <= 8'h87;
			14'd11438: ff_rdata <= 8'h87;
			14'd11439: ff_rdata <= 8'h67;
			14'd11440: ff_rdata <= 8'h87;
			14'd11441: ff_rdata <= 8'h84;
			14'd11442: ff_rdata <= 8'h21;
			14'd11443: ff_rdata <= 8'hD2;
			14'd11444: ff_rdata <= 8'h6C;
			14'd11445: ff_rdata <= 8'hCD;
			14'd11446: ff_rdata <= 8'h86;
			14'd11447: ff_rdata <= 8'h54;
			14'd11448: ff_rdata <= 8'h11;
			14'd11449: ff_rdata <= 8'h09;
			14'd11450: ff_rdata <= 8'h00;
			14'd11451: ff_rdata <= 8'h19;
			14'd11452: ff_rdata <= 8'h4E;
			14'd11453: ff_rdata <= 8'hED;
			14'd11454: ff_rdata <= 8'h52;
			14'd11455: ff_rdata <= 8'h11;
			14'd11456: ff_rdata <= 8'hA3;
			14'd11457: ff_rdata <= 8'hF9;
			14'd11458: ff_rdata <= 8'hED;
			14'd11459: ff_rdata <= 8'h53;
			14'd11460: ff_rdata <= 8'hA1;
			14'd11461: ff_rdata <= 8'hF9;
			14'd11462: ff_rdata <= 8'h06;
			14'd11463: ff_rdata <= 8'h0C;
			14'd11464: ff_rdata <= 8'h7E;
			14'd11465: ff_rdata <= 8'h91;
			14'd11466: ff_rdata <= 8'h12;
			14'd11467: ff_rdata <= 8'h23;
			14'd11468: ff_rdata <= 8'h13;
			14'd11469: ff_rdata <= 8'h10;
			14'd11470: ff_rdata <= 8'hF9;
			14'd11471: ff_rdata <= 8'hE1;
			14'd11472: ff_rdata <= 8'hA7;
			14'd11473: ff_rdata <= 8'hC9;
			14'd11474: ff_rdata <= 8'hF1;
			14'd11475: ff_rdata <= 8'h14;
			14'd11476: ff_rdata <= 8'hFB;
			14'd11477: ff_rdata <= 8'hE2;
			14'd11478: ff_rdata <= 8'h05;
			14'd11479: ff_rdata <= 8'hEC;
			14'd11480: ff_rdata <= 8'h0F;
			14'd11481: ff_rdata <= 8'hF6;
			14'd11482: ff_rdata <= 8'h19;
			14'd11483: ff_rdata <= 8'h00;
			14'd11484: ff_rdata <= 8'hE7;
			14'd11485: ff_rdata <= 8'h0A;
			14'd11486: ff_rdata <= 8'h1A;
			14'd11487: ff_rdata <= 8'hDD;
			14'd11488: ff_rdata <= 8'h09;
			14'd11489: ff_rdata <= 8'h35;
			14'd11490: ff_rdata <= 8'hF7;
			14'd11491: ff_rdata <= 8'h23;
			14'd11492: ff_rdata <= 8'hE6;
			14'd11493: ff_rdata <= 8'h12;
			14'd11494: ff_rdata <= 8'hD4;
			14'd11495: ff_rdata <= 8'h00;
			14'd11496: ff_rdata <= 8'h2C;
			14'd11497: ff_rdata <= 8'hEE;
			14'd11498: ff_rdata <= 8'h1E;
			14'd11499: ff_rdata <= 8'h05;
			14'd11500: ff_rdata <= 8'h0A;
			14'd11501: ff_rdata <= 8'h0F;
			14'd11502: ff_rdata <= 8'h05;
			14'd11503: ff_rdata <= 8'h19;
			14'd11504: ff_rdata <= 8'h00;
			14'd11505: ff_rdata <= 8'h14;
			14'd11506: ff_rdata <= 8'h0A;
			14'd11507: ff_rdata <= 8'h00;
			14'd11508: ff_rdata <= 8'h14;
			14'd11509: ff_rdata <= 8'h0A;
			14'd11510: ff_rdata <= 8'h1E;
			14'd11511: ff_rdata <= 8'h05;
			14'd11512: ff_rdata <= 8'h0A;
			14'd11513: ff_rdata <= 8'h0F;
			14'd11514: ff_rdata <= 8'h05;
			14'd11515: ff_rdata <= 8'h19;
			14'd11516: ff_rdata <= 8'h00;
			14'd11517: ff_rdata <= 8'h14;
			14'd11518: ff_rdata <= 8'h0A;
			14'd11519: ff_rdata <= 8'h00;
			14'd11520: ff_rdata <= 8'h14;
			14'd11521: ff_rdata <= 8'hFB;
			14'd11522: ff_rdata <= 8'h00;
			14'd11523: ff_rdata <= 8'hF6;
			14'd11524: ff_rdata <= 8'h0A;
			14'd11525: ff_rdata <= 8'h00;
			14'd11526: ff_rdata <= 8'hF6;
			14'd11527: ff_rdata <= 8'h0A;
			14'd11528: ff_rdata <= 8'h00;
			14'd11529: ff_rdata <= 8'h05;
			14'd11530: ff_rdata <= 8'hEC;
			14'd11531: ff_rdata <= 8'h00;
			14'd11532: ff_rdata <= 8'h05;
			14'd11533: ff_rdata <= 8'hFB;
			14'd11534: ff_rdata <= 8'h1A;
			14'd11535: ff_rdata <= 8'h01;
			14'd11536: ff_rdata <= 8'h09;
			14'd11537: ff_rdata <= 8'h0B;
			14'd11538: ff_rdata <= 8'hF7;
			14'd11539: ff_rdata <= 8'h15;
			14'd11540: ff_rdata <= 8'h01;
			14'd11541: ff_rdata <= 8'h12;
			14'd11542: ff_rdata <= 8'h06;
			14'd11543: ff_rdata <= 8'h00;
			14'd11544: ff_rdata <= 8'h10;
			14'd11545: ff_rdata <= 8'hFC;
			14'd11546: ff_rdata <= 8'h1A;
			14'd11547: ff_rdata <= 8'h01;
			14'd11548: ff_rdata <= 8'h09;
			14'd11549: ff_rdata <= 8'h0B;
			14'd11550: ff_rdata <= 8'h05;
			14'd11551: ff_rdata <= 8'h15;
			14'd11552: ff_rdata <= 8'h01;
			14'd11553: ff_rdata <= 8'h12;
			14'd11554: ff_rdata <= 8'h06;
			14'd11555: ff_rdata <= 8'h00;
			14'd11556: ff_rdata <= 8'h10;
			14'd11557: ff_rdata <= 8'h0A;
			14'd11558: ff_rdata <= 8'h0F;
			14'd11559: ff_rdata <= 8'h00;
			14'd11560: ff_rdata <= 8'h05;
			14'd11561: ff_rdata <= 8'h0A;
			14'd11562: ff_rdata <= 8'hFB;
			14'd11563: ff_rdata <= 8'h14;
			14'd11564: ff_rdata <= 8'hFB;
			14'd11565: ff_rdata <= 8'h0A;
			14'd11566: ff_rdata <= 8'h05;
			14'd11567: ff_rdata <= 8'h00;
			14'd11568: ff_rdata <= 8'h0F;
			14'd11569: ff_rdata <= 8'hF6;
			14'd11570: ff_rdata <= 8'h1A;
			14'd11571: ff_rdata <= 8'hF8;
			14'd11572: ff_rdata <= 8'h09;
			14'd11573: ff_rdata <= 8'h27;
			14'd11574: ff_rdata <= 8'hF7;
			14'd11575: ff_rdata <= 8'h23;
			14'd11576: ff_rdata <= 8'hF3;
			14'd11577: ff_rdata <= 8'h12;
			14'd11578: ff_rdata <= 8'hFD;
			14'd11579: ff_rdata <= 8'h00;
			14'd11580: ff_rdata <= 8'h2C;
			14'd11581: ff_rdata <= 8'hEE;
			14'd11582: ff_rdata <= 8'h00;
			14'd11583: ff_rdata <= 8'h00;
			14'd11584: ff_rdata <= 8'h00;
			14'd11585: ff_rdata <= 8'h00;
			14'd11586: ff_rdata <= 8'h00;
			14'd11587: ff_rdata <= 8'h00;
			14'd11588: ff_rdata <= 8'h00;
			14'd11589: ff_rdata <= 8'h00;
			14'd11590: ff_rdata <= 8'h00;
			14'd11591: ff_rdata <= 8'h00;
			14'd11592: ff_rdata <= 8'h00;
			14'd11593: ff_rdata <= 8'h00;
			14'd11594: ff_rdata <= 8'h29;
			14'd11595: ff_rdata <= 8'hDC;
			14'd11596: ff_rdata <= 8'h33;
			14'd11597: ff_rdata <= 8'h52;
			14'd11598: ff_rdata <= 8'h05;
			14'd11599: ff_rdata <= 8'h24;
			14'd11600: ff_rdata <= 8'hD7;
			14'd11601: ff_rdata <= 8'h2E;
			14'd11602: ff_rdata <= 8'hE1;
			14'd11603: ff_rdata <= 8'h00;
			14'd11604: ff_rdata <= 8'h56;
			14'd11605: ff_rdata <= 8'h0A;
			14'd11606: ff_rdata <= 8'h29;
			14'd11607: ff_rdata <= 8'hDC;
			14'd11608: ff_rdata <= 8'h33;
			14'd11609: ff_rdata <= 8'h52;
			14'd11610: ff_rdata <= 8'h05;
			14'd11611: ff_rdata <= 8'h24;
			14'd11612: ff_rdata <= 8'hD7;
			14'd11613: ff_rdata <= 8'h2E;
			14'd11614: ff_rdata <= 8'hE1;
			14'd11615: ff_rdata <= 8'h00;
			14'd11616: ff_rdata <= 8'h56;
			14'd11617: ff_rdata <= 8'hAF;
			14'd11618: ff_rdata <= 8'h0E;
			14'd11619: ff_rdata <= 8'h00;
			14'd11620: ff_rdata <= 8'h06;
			14'd11621: ff_rdata <= 8'h08;
			14'd11622: ff_rdata <= 8'hCD;
			14'd11623: ff_rdata <= 8'h7B;
			14'd11624: ff_rdata <= 8'h6D;
			14'd11625: ff_rdata <= 8'h0E;
			14'd11626: ff_rdata <= 8'h0E;
			14'd11627: ff_rdata <= 8'h06;
			14'd11628: ff_rdata <= 8'h0B;
			14'd11629: ff_rdata <= 8'hCD;
			14'd11630: ff_rdata <= 8'h7B;
			14'd11631: ff_rdata <= 8'h6D;
			14'd11632: ff_rdata <= 8'h0E;
			14'd11633: ff_rdata <= 8'h20;
			14'd11634: ff_rdata <= 8'h06;
			14'd11635: ff_rdata <= 8'h09;
			14'd11636: ff_rdata <= 8'hCD;
			14'd11637: ff_rdata <= 8'h7B;
			14'd11638: ff_rdata <= 8'h6D;
			14'd11639: ff_rdata <= 8'h0E;
			14'd11640: ff_rdata <= 8'h30;
			14'd11641: ff_rdata <= 8'h06;
			14'd11642: ff_rdata <= 8'h09;
			14'd11643: ff_rdata <= 8'hC5;
			14'd11644: ff_rdata <= 8'h47;
			14'd11645: ff_rdata <= 8'hCD;
			14'd11646: ff_rdata <= 8'hB5;
			14'd11647: ff_rdata <= 8'h6D;
			14'd11648: ff_rdata <= 8'hFB;
			14'd11649: ff_rdata <= 8'hC1;
			14'd11650: ff_rdata <= 8'h0C;
			14'd11651: ff_rdata <= 8'h10;
			14'd11652: ff_rdata <= 8'hF6;
			14'd11653: ff_rdata <= 8'hC9;
			14'd11654: ff_rdata <= 8'h0E;
			14'd11655: ff_rdata <= 8'h0E;
			14'd11656: ff_rdata <= 8'hCD;
			14'd11657: ff_rdata <= 8'hE0;
			14'd11658: ff_rdata <= 8'h6D;
			14'd11659: ff_rdata <= 8'hF6;
			14'd11660: ff_rdata <= 8'h20;
			14'd11661: ff_rdata <= 8'h47;
			14'd11662: ff_rdata <= 8'hCD;
			14'd11663: ff_rdata <= 8'hB5;
			14'd11664: ff_rdata <= 8'h6D;
			14'd11665: ff_rdata <= 8'h21;
			14'd11666: ff_rdata <= 8'hA3;
			14'd11667: ff_rdata <= 8'h6D;
			14'd11668: ff_rdata <= 8'h06;
			14'd11669: ff_rdata <= 8'h09;
			14'd11670: ff_rdata <= 8'hC5;
			14'd11671: ff_rdata <= 8'h4E;
			14'd11672: ff_rdata <= 8'h23;
			14'd11673: ff_rdata <= 8'h46;
			14'd11674: ff_rdata <= 8'h23;
			14'd11675: ff_rdata <= 8'hCD;
			14'd11676: ff_rdata <= 8'hB5;
			14'd11677: ff_rdata <= 8'h6D;
			14'd11678: ff_rdata <= 8'hFB;
			14'd11679: ff_rdata <= 8'hC1;
			14'd11680: ff_rdata <= 8'h10;
			14'd11681: ff_rdata <= 8'hF4;
			14'd11682: ff_rdata <= 8'hC9;
			14'd11683: ff_rdata <= 8'h16;
			14'd11684: ff_rdata <= 8'h20;
			14'd11685: ff_rdata <= 8'h17;
			14'd11686: ff_rdata <= 8'h50;
			14'd11687: ff_rdata <= 8'h18;
			14'd11688: ff_rdata <= 8'hC0;
			14'd11689: ff_rdata <= 8'h26;
			14'd11690: ff_rdata <= 8'h05;
			14'd11691: ff_rdata <= 8'h27;
			14'd11692: ff_rdata <= 8'h05;
			14'd11693: ff_rdata <= 8'h28;
			14'd11694: ff_rdata <= 8'h01;
			14'd11695: ff_rdata <= 8'h36;
			14'd11696: ff_rdata <= 8'h00;
			14'd11697: ff_rdata <= 8'h37;
			14'd11698: ff_rdata <= 8'h00;
			14'd11699: ff_rdata <= 8'h38;
			14'd11700: ff_rdata <= 8'h00;
			14'd11701: ff_rdata <= 8'hF5;
			14'd11702: ff_rdata <= 8'h79;
			14'd11703: ff_rdata <= 8'hCD;
			14'd11704: ff_rdata <= 8'hF3;
			14'd11705: ff_rdata <= 8'h6D;
			14'd11706: ff_rdata <= 8'h38;
			14'd11707: ff_rdata <= 8'h21;
			14'd11708: ff_rdata <= 8'hE5;
			14'd11709: ff_rdata <= 8'h21;
			14'd11710: ff_rdata <= 8'hC0;
			14'd11711: ff_rdata <= 8'hF9;
			14'd11712: ff_rdata <= 8'h85;
			14'd11713: ff_rdata <= 8'h6F;
			14'd11714: ff_rdata <= 8'h3E;
			14'd11715: ff_rdata <= 8'h00;
			14'd11716: ff_rdata <= 8'h8C;
			14'd11717: ff_rdata <= 8'h67;
			14'd11718: ff_rdata <= 8'hF3;
			14'd11719: ff_rdata <= 8'h70;
			14'd11720: ff_rdata <= 8'h79;
			14'd11721: ff_rdata <= 8'hD3;
			14'd11722: ff_rdata <= 8'h7C;
			14'd11723: ff_rdata <= 8'hE3;
			14'd11724: ff_rdata <= 8'hE3;
			14'd11725: ff_rdata <= 8'h78;
			14'd11726: ff_rdata <= 8'hD3;
			14'd11727: ff_rdata <= 8'h7D;
			14'd11728: ff_rdata <= 8'hE3;
			14'd11729: ff_rdata <= 8'hE3;
			14'd11730: ff_rdata <= 8'hE3;
			14'd11731: ff_rdata <= 8'hE3;
			14'd11732: ff_rdata <= 8'hE3;
			14'd11733: ff_rdata <= 8'hE3;
			14'd11734: ff_rdata <= 8'hE3;
			14'd11735: ff_rdata <= 8'hE3;
			14'd11736: ff_rdata <= 8'hE1;
			14'd11737: ff_rdata <= 8'hF1;
			14'd11738: ff_rdata <= 8'h37;
			14'd11739: ff_rdata <= 8'h3F;
			14'd11740: ff_rdata <= 8'hC9;
			14'd11741: ff_rdata <= 8'hF1;
			14'd11742: ff_rdata <= 8'h37;
			14'd11743: ff_rdata <= 8'hC9;
			14'd11744: ff_rdata <= 8'h79;
			14'd11745: ff_rdata <= 8'hCD;
			14'd11746: ff_rdata <= 8'hF3;
			14'd11747: ff_rdata <= 8'h6D;
			14'd11748: ff_rdata <= 8'hD8;
			14'd11749: ff_rdata <= 8'hE5;
			14'd11750: ff_rdata <= 8'h21;
			14'd11751: ff_rdata <= 8'hC0;
			14'd11752: ff_rdata <= 8'hF9;
			14'd11753: ff_rdata <= 8'h79;
			14'd11754: ff_rdata <= 8'h85;
			14'd11755: ff_rdata <= 8'h6F;
			14'd11756: ff_rdata <= 8'h3E;
			14'd11757: ff_rdata <= 8'h00;
			14'd11758: ff_rdata <= 8'h8C;
			14'd11759: ff_rdata <= 8'h67;
			14'd11760: ff_rdata <= 8'h7E;
			14'd11761: ff_rdata <= 8'hE1;
			14'd11762: ff_rdata <= 8'hC9;
			14'd11763: ff_rdata <= 8'hFE;
			14'd11764: ff_rdata <= 8'h08;
			14'd11765: ff_rdata <= 8'h3F;
			14'd11766: ff_rdata <= 8'hD0;
			14'd11767: ff_rdata <= 8'hFE;
			14'd11768: ff_rdata <= 8'h0E;
			14'd11769: ff_rdata <= 8'hD8;
			14'd11770: ff_rdata <= 8'hFE;
			14'd11771: ff_rdata <= 8'h19;
			14'd11772: ff_rdata <= 8'h3F;
			14'd11773: ff_rdata <= 8'hD0;
			14'd11774: ff_rdata <= 8'hFE;
			14'd11775: ff_rdata <= 8'h20;
			14'd11776: ff_rdata <= 8'hD8;
			14'd11777: ff_rdata <= 8'hFE;
			14'd11778: ff_rdata <= 8'h29;
			14'd11779: ff_rdata <= 8'h3F;
			14'd11780: ff_rdata <= 8'hD0;
			14'd11781: ff_rdata <= 8'hFE;
			14'd11782: ff_rdata <= 8'h30;
			14'd11783: ff_rdata <= 8'hD8;
			14'd11784: ff_rdata <= 8'hFE;
			14'd11785: ff_rdata <= 8'h39;
			14'd11786: ff_rdata <= 8'h3F;
			14'd11787: ff_rdata <= 8'hC9;
			14'd11788: ff_rdata <= 8'h50;
			14'd11789: ff_rdata <= 8'h69;
			14'd11790: ff_rdata <= 8'h61;
			14'd11791: ff_rdata <= 8'h6E;
			14'd11792: ff_rdata <= 8'h6F;
			14'd11793: ff_rdata <= 8'h20;
			14'd11794: ff_rdata <= 8'h31;
			14'd11795: ff_rdata <= 8'h20;
			14'd11796: ff_rdata <= 8'h00;
			14'd11797: ff_rdata <= 8'h00;
			14'd11798: ff_rdata <= 8'h0A;
			14'd11799: ff_rdata <= 8'h00;
			14'd11800: ff_rdata <= 8'h00;
			14'd11801: ff_rdata <= 8'h00;
			14'd11802: ff_rdata <= 8'h00;
			14'd11803: ff_rdata <= 8'h00;
			14'd11804: ff_rdata <= 8'h31;
			14'd11805: ff_rdata <= 8'h0E;
			14'd11806: ff_rdata <= 8'hD9;
			14'd11807: ff_rdata <= 8'h11;
			14'd11808: ff_rdata <= 8'h30;
			14'd11809: ff_rdata <= 8'h00;
			14'd11810: ff_rdata <= 8'h00;
			14'd11811: ff_rdata <= 8'h00;
			14'd11812: ff_rdata <= 8'h11;
			14'd11813: ff_rdata <= 8'h00;
			14'd11814: ff_rdata <= 8'hB2;
			14'd11815: ff_rdata <= 8'hF4;
			14'd11816: ff_rdata <= 8'h70;
			14'd11817: ff_rdata <= 8'h00;
			14'd11818: ff_rdata <= 8'h00;
			14'd11819: ff_rdata <= 8'h00;
			14'd11820: ff_rdata <= 8'h50;
			14'd11821: ff_rdata <= 8'h69;
			14'd11822: ff_rdata <= 8'h61;
			14'd11823: ff_rdata <= 8'h6E;
			14'd11824: ff_rdata <= 8'h6F;
			14'd11825: ff_rdata <= 8'h20;
			14'd11826: ff_rdata <= 8'h32;
			14'd11827: ff_rdata <= 8'h20;
			14'd11828: ff_rdata <= 8'h00;
			14'd11829: ff_rdata <= 8'h0C;
			14'd11830: ff_rdata <= 8'h08;
			14'd11831: ff_rdata <= 8'h00;
			14'd11832: ff_rdata <= 8'h00;
			14'd11833: ff_rdata <= 8'h00;
			14'd11834: ff_rdata <= 8'h00;
			14'd11835: ff_rdata <= 8'h00;
			14'd11836: ff_rdata <= 8'h30;
			14'd11837: ff_rdata <= 8'h0F;
			14'd11838: ff_rdata <= 8'hD9;
			14'd11839: ff_rdata <= 8'h10;
			14'd11840: ff_rdata <= 8'h30;
			14'd11841: ff_rdata <= 8'h00;
			14'd11842: ff_rdata <= 8'h00;
			14'd11843: ff_rdata <= 8'h00;
			14'd11844: ff_rdata <= 8'h10;
			14'd11845: ff_rdata <= 8'h00;
			14'd11846: ff_rdata <= 8'hB2;
			14'd11847: ff_rdata <= 8'hF3;
			14'd11848: ff_rdata <= 8'h70;
			14'd11849: ff_rdata <= 8'h00;
			14'd11850: ff_rdata <= 8'h00;
			14'd11851: ff_rdata <= 8'h00;
			14'd11852: ff_rdata <= 8'h56;
			14'd11853: ff_rdata <= 8'h69;
			14'd11854: ff_rdata <= 8'h6F;
			14'd11855: ff_rdata <= 8'h6C;
			14'd11856: ff_rdata <= 8'h69;
			14'd11857: ff_rdata <= 8'h6E;
			14'd11858: ff_rdata <= 8'h20;
			14'd11859: ff_rdata <= 8'h20;
			14'd11860: ff_rdata <= 8'h00;
			14'd11861: ff_rdata <= 8'h0C;
			14'd11862: ff_rdata <= 8'h6E;
			14'd11863: ff_rdata <= 8'h00;
			14'd11864: ff_rdata <= 8'h00;
			14'd11865: ff_rdata <= 8'h00;
			14'd11866: ff_rdata <= 8'h00;
			14'd11867: ff_rdata <= 8'h00;
			14'd11868: ff_rdata <= 8'h61;
			14'd11869: ff_rdata <= 8'h12;
			14'd11870: ff_rdata <= 8'hB4;
			14'd11871: ff_rdata <= 8'h14;
			14'd11872: ff_rdata <= 8'h10;
			14'd11873: ff_rdata <= 8'h00;
			14'd11874: ff_rdata <= 8'h00;
			14'd11875: ff_rdata <= 8'h00;
			14'd11876: ff_rdata <= 8'h61;
			14'd11877: ff_rdata <= 8'h00;
			14'd11878: ff_rdata <= 8'h56;
			14'd11879: ff_rdata <= 8'h17;
			14'd11880: ff_rdata <= 8'h80;
			14'd11881: ff_rdata <= 8'h00;
			14'd11882: ff_rdata <= 8'h00;
			14'd11883: ff_rdata <= 8'h00;
			14'd11884: ff_rdata <= 8'h46;
			14'd11885: ff_rdata <= 8'h6C;
			14'd11886: ff_rdata <= 8'h75;
			14'd11887: ff_rdata <= 8'h74;
			14'd11888: ff_rdata <= 8'h65;
			14'd11889: ff_rdata <= 8'h20;
			14'd11890: ff_rdata <= 8'h20;
			14'd11891: ff_rdata <= 8'h20;
			14'd11892: ff_rdata <= 8'h00;
			14'd11893: ff_rdata <= 8'h0C;
			14'd11894: ff_rdata <= 8'h0E;
			14'd11895: ff_rdata <= 8'h00;
			14'd11896: ff_rdata <= 8'h00;
			14'd11897: ff_rdata <= 8'h00;
			14'd11898: ff_rdata <= 8'h00;
			14'd11899: ff_rdata <= 8'h00;
			14'd11900: ff_rdata <= 8'h61;
			14'd11901: ff_rdata <= 8'h20;
			14'd11902: ff_rdata <= 8'h6C;
			14'd11903: ff_rdata <= 8'h18;
			14'd11904: ff_rdata <= 8'h40;
			14'd11905: ff_rdata <= 8'h00;
			14'd11906: ff_rdata <= 8'h00;
			14'd11907: ff_rdata <= 8'h00;
			14'd11908: ff_rdata <= 8'h31;
			14'd11909: ff_rdata <= 8'h03;
			14'd11910: ff_rdata <= 8'h43;
			14'd11911: ff_rdata <= 8'h26;
			14'd11912: ff_rdata <= 8'h80;
			14'd11913: ff_rdata <= 8'h00;
			14'd11914: ff_rdata <= 8'h00;
			14'd11915: ff_rdata <= 8'h00;
			14'd11916: ff_rdata <= 8'h43;
			14'd11917: ff_rdata <= 8'h6C;
			14'd11918: ff_rdata <= 8'h61;
			14'd11919: ff_rdata <= 8'h72;
			14'd11920: ff_rdata <= 8'h69;
			14'd11921: ff_rdata <= 8'h6E;
			14'd11922: ff_rdata <= 8'h65;
			14'd11923: ff_rdata <= 8'h74;
			14'd11924: ff_rdata <= 8'h00;
			14'd11925: ff_rdata <= 8'h0C;
			14'd11926: ff_rdata <= 8'h0E;
			14'd11927: ff_rdata <= 8'h00;
			14'd11928: ff_rdata <= 8'h00;
			14'd11929: ff_rdata <= 8'h00;
			14'd11930: ff_rdata <= 8'h00;
			14'd11931: ff_rdata <= 8'h00;
			14'd11932: ff_rdata <= 8'hA2;
			14'd11933: ff_rdata <= 8'hA0;
			14'd11934: ff_rdata <= 8'h88;
			14'd11935: ff_rdata <= 8'h14;
			14'd11936: ff_rdata <= 8'h40;
			14'd11937: ff_rdata <= 8'h00;
			14'd11938: ff_rdata <= 8'h00;
			14'd11939: ff_rdata <= 8'h00;
			14'd11940: ff_rdata <= 8'h30;
			14'd11941: ff_rdata <= 8'h00;
			14'd11942: ff_rdata <= 8'h54;
			14'd11943: ff_rdata <= 8'h06;
			14'd11944: ff_rdata <= 8'h80;
			14'd11945: ff_rdata <= 8'h00;
			14'd11946: ff_rdata <= 8'h00;
			14'd11947: ff_rdata <= 8'h00;
			14'd11948: ff_rdata <= 8'h4F;
			14'd11949: ff_rdata <= 8'h62;
			14'd11950: ff_rdata <= 8'h6F;
			14'd11951: ff_rdata <= 8'h65;
			14'd11952: ff_rdata <= 8'h20;
			14'd11953: ff_rdata <= 8'h20;
			14'd11954: ff_rdata <= 8'h20;
			14'd11955: ff_rdata <= 8'h20;
			14'd11956: ff_rdata <= 8'h00;
			14'd11957: ff_rdata <= 8'h00;
			14'd11958: ff_rdata <= 8'h0A;
			14'd11959: ff_rdata <= 8'h00;
			14'd11960: ff_rdata <= 8'h00;
			14'd11961: ff_rdata <= 8'h00;
			14'd11962: ff_rdata <= 8'h00;
			14'd11963: ff_rdata <= 8'h00;
			14'd11964: ff_rdata <= 8'h31;
			14'd11965: ff_rdata <= 8'h20;
			14'd11966: ff_rdata <= 8'h72;
			14'd11967: ff_rdata <= 8'h0A;
			14'd11968: ff_rdata <= 8'h40;
			14'd11969: ff_rdata <= 8'h00;
			14'd11970: ff_rdata <= 8'h00;
			14'd11971: ff_rdata <= 8'h00;
			14'd11972: ff_rdata <= 8'h34;
			14'd11973: ff_rdata <= 8'h01;
			14'd11974: ff_rdata <= 8'h56;
			14'd11975: ff_rdata <= 8'h1C;
			14'd11976: ff_rdata <= 8'h80;
			14'd11977: ff_rdata <= 8'h00;
			14'd11978: ff_rdata <= 8'h00;
			14'd11979: ff_rdata <= 8'h00;
			14'd11980: ff_rdata <= 8'h54;
			14'd11981: ff_rdata <= 8'h72;
			14'd11982: ff_rdata <= 8'h75;
			14'd11983: ff_rdata <= 8'h6D;
			14'd11984: ff_rdata <= 8'h70;
			14'd11985: ff_rdata <= 8'h65;
			14'd11986: ff_rdata <= 8'h74;
			14'd11987: ff_rdata <= 8'h20;
			14'd11988: ff_rdata <= 8'h00;
			14'd11989: ff_rdata <= 8'h00;
			14'd11990: ff_rdata <= 8'h6E;
			14'd11991: ff_rdata <= 8'h00;
			14'd11992: ff_rdata <= 8'h00;
			14'd11993: ff_rdata <= 8'h00;
			14'd11994: ff_rdata <= 8'h00;
			14'd11995: ff_rdata <= 8'h00;
			14'd11996: ff_rdata <= 8'h31;
			14'd11997: ff_rdata <= 8'h16;
			14'd11998: ff_rdata <= 8'h51;
			14'd11999: ff_rdata <= 8'h26;
			14'd12000: ff_rdata <= 8'h40;
			14'd12001: ff_rdata <= 8'h00;
			14'd12002: ff_rdata <= 8'h00;
			14'd12003: ff_rdata <= 8'h00;
			14'd12004: ff_rdata <= 8'h71;
			14'd12005: ff_rdata <= 8'h03;
			14'd12006: ff_rdata <= 8'h52;
			14'd12007: ff_rdata <= 8'h24;
			14'd12008: ff_rdata <= 8'h60;
			14'd12009: ff_rdata <= 8'h00;
			14'd12010: ff_rdata <= 8'h00;
			14'd12011: ff_rdata <= 8'h00;
			14'd12012: ff_rdata <= 8'h50;
			14'd12013: ff_rdata <= 8'h69;
			14'd12014: ff_rdata <= 8'h70;
			14'd12015: ff_rdata <= 8'h65;
			14'd12016: ff_rdata <= 8'h4F;
			14'd12017: ff_rdata <= 8'h72;
			14'd12018: ff_rdata <= 8'h67;
			14'd12019: ff_rdata <= 8'h6E;
			14'd12020: ff_rdata <= 8'h01;
			14'd12021: ff_rdata <= 8'h00;
			14'd12022: ff_rdata <= 8'h0C;
			14'd12023: ff_rdata <= 8'h00;
			14'd12024: ff_rdata <= 8'h00;
			14'd12025: ff_rdata <= 8'h00;
			14'd12026: ff_rdata <= 8'h00;
			14'd12027: ff_rdata <= 8'h00;
			14'd12028: ff_rdata <= 8'h34;
			14'd12029: ff_rdata <= 8'h37;
			14'd12030: ff_rdata <= 8'h50;
			14'd12031: ff_rdata <= 8'h76;
			14'd12032: ff_rdata <= 8'h30;
			14'd12033: ff_rdata <= 8'h00;
			14'd12034: ff_rdata <= 8'h00;
			14'd12035: ff_rdata <= 8'h00;
			14'd12036: ff_rdata <= 8'h30;
			14'd12037: ff_rdata <= 8'h00;
			14'd12038: ff_rdata <= 8'h30;
			14'd12039: ff_rdata <= 8'h06;
			14'd12040: ff_rdata <= 8'h80;
			14'd12041: ff_rdata <= 8'h00;
			14'd12042: ff_rdata <= 8'h00;
			14'd12043: ff_rdata <= 8'h00;
			14'd12044: ff_rdata <= 8'h58;
			14'd12045: ff_rdata <= 8'h79;
			14'd12046: ff_rdata <= 8'h6C;
			14'd12047: ff_rdata <= 8'h6F;
			14'd12048: ff_rdata <= 8'h70;
			14'd12049: ff_rdata <= 8'h68;
			14'd12050: ff_rdata <= 8'h6F;
			14'd12051: ff_rdata <= 8'h6E;
			14'd12052: ff_rdata <= 8'h00;
			14'd12053: ff_rdata <= 8'h00;
			14'd12054: ff_rdata <= 8'h0A;
			14'd12055: ff_rdata <= 8'h00;
			14'd12056: ff_rdata <= 8'h00;
			14'd12057: ff_rdata <= 8'h00;
			14'd12058: ff_rdata <= 8'h00;
			14'd12059: ff_rdata <= 8'h00;
			14'd12060: ff_rdata <= 8'h17;
			14'd12061: ff_rdata <= 8'h18;
			14'd12062: ff_rdata <= 8'h88;
			14'd12063: ff_rdata <= 8'h66;
			14'd12064: ff_rdata <= 8'h80;
			14'd12065: ff_rdata <= 8'h00;
			14'd12066: ff_rdata <= 8'h00;
			14'd12067: ff_rdata <= 8'h00;
			14'd12068: ff_rdata <= 8'h52;
			14'd12069: ff_rdata <= 8'h00;
			14'd12070: ff_rdata <= 8'hD9;
			14'd12071: ff_rdata <= 8'h24;
			14'd12072: ff_rdata <= 8'h80;
			14'd12073: ff_rdata <= 8'h00;
			14'd12074: ff_rdata <= 8'h00;
			14'd12075: ff_rdata <= 8'h00;
			14'd12076: ff_rdata <= 8'h4F;
			14'd12077: ff_rdata <= 8'h72;
			14'd12078: ff_rdata <= 8'h67;
			14'd12079: ff_rdata <= 8'h61;
			14'd12080: ff_rdata <= 8'h6E;
			14'd12081: ff_rdata <= 8'h20;
			14'd12082: ff_rdata <= 8'h20;
			14'd12083: ff_rdata <= 8'h20;
			14'd12084: ff_rdata <= 8'h00;
			14'd12085: ff_rdata <= 8'h00;
			14'd12086: ff_rdata <= 8'hED;
			14'd12087: ff_rdata <= 8'h00;
			14'd12088: ff_rdata <= 8'h00;
			14'd12089: ff_rdata <= 8'h00;
			14'd12090: ff_rdata <= 8'h00;
			14'd12091: ff_rdata <= 8'h00;
			14'd12092: ff_rdata <= 8'hE1;
			14'd12093: ff_rdata <= 8'h0A;
			14'd12094: ff_rdata <= 8'hFC;
			14'd12095: ff_rdata <= 8'h28;
			14'd12096: ff_rdata <= 8'h70;
			14'd12097: ff_rdata <= 8'h00;
			14'd12098: ff_rdata <= 8'h00;
			14'd12099: ff_rdata <= 8'h00;
			14'd12100: ff_rdata <= 8'h63;
			14'd12101: ff_rdata <= 8'h05;
			14'd12102: ff_rdata <= 8'hF8;
			14'd12103: ff_rdata <= 8'h29;
			14'd12104: ff_rdata <= 8'h70;
			14'd12105: ff_rdata <= 8'h00;
			14'd12106: ff_rdata <= 8'h00;
			14'd12107: ff_rdata <= 8'h00;
			14'd12108: ff_rdata <= 8'h47;
			14'd12109: ff_rdata <= 8'h75;
			14'd12110: ff_rdata <= 8'h69;
			14'd12111: ff_rdata <= 8'h74;
			14'd12112: ff_rdata <= 8'h61;
			14'd12113: ff_rdata <= 8'h72;
			14'd12114: ff_rdata <= 8'h20;
			14'd12115: ff_rdata <= 8'h20;
			14'd12116: ff_rdata <= 8'h00;
			14'd12117: ff_rdata <= 8'h00;
			14'd12118: ff_rdata <= 8'h0A;
			14'd12119: ff_rdata <= 8'h00;
			14'd12120: ff_rdata <= 8'h00;
			14'd12121: ff_rdata <= 8'h00;
			14'd12122: ff_rdata <= 8'h00;
			14'd12123: ff_rdata <= 8'h00;
			14'd12124: ff_rdata <= 8'h02;
			14'd12125: ff_rdata <= 8'h15;
			14'd12126: ff_rdata <= 8'hA3;
			14'd12127: ff_rdata <= 8'h75;
			14'd12128: ff_rdata <= 8'h20;
			14'd12129: ff_rdata <= 8'h00;
			14'd12130: ff_rdata <= 8'h00;
			14'd12131: ff_rdata <= 8'h00;
			14'd12132: ff_rdata <= 8'h41;
			14'd12133: ff_rdata <= 8'h00;
			14'd12134: ff_rdata <= 8'hA3;
			14'd12135: ff_rdata <= 8'h05;
			14'd12136: ff_rdata <= 8'h60;
			14'd12137: ff_rdata <= 8'h00;
			14'd12138: ff_rdata <= 8'h00;
			14'd12139: ff_rdata <= 8'h00;
			14'd12140: ff_rdata <= 8'h53;
			14'd12141: ff_rdata <= 8'h61;
			14'd12142: ff_rdata <= 8'h6E;
			14'd12143: ff_rdata <= 8'h74;
			14'd12144: ff_rdata <= 8'h6F;
			14'd12145: ff_rdata <= 8'h6F;
			14'd12146: ff_rdata <= 8'h6C;
			14'd12147: ff_rdata <= 8'h20;
			14'd12148: ff_rdata <= 8'h00;
			14'd12149: ff_rdata <= 8'hF9;
			14'd12150: ff_rdata <= 8'h0C;
			14'd12151: ff_rdata <= 8'h00;
			14'd12152: ff_rdata <= 8'h00;
			14'd12153: ff_rdata <= 8'h00;
			14'd12154: ff_rdata <= 8'h00;
			14'd12155: ff_rdata <= 8'h00;
			14'd12156: ff_rdata <= 8'h19;
			14'd12157: ff_rdata <= 8'h0C;
			14'd12158: ff_rdata <= 8'hC7;
			14'd12159: ff_rdata <= 8'h11;
			14'd12160: ff_rdata <= 8'h10;
			14'd12161: ff_rdata <= 8'h00;
			14'd12162: ff_rdata <= 8'h00;
			14'd12163: ff_rdata <= 8'h00;
			14'd12164: ff_rdata <= 8'h53;
			14'd12165: ff_rdata <= 8'h03;
			14'd12166: ff_rdata <= 8'hF5;
			14'd12167: ff_rdata <= 8'h03;
			14'd12168: ff_rdata <= 8'h60;
			14'd12169: ff_rdata <= 8'h00;
			14'd12170: ff_rdata <= 8'h00;
			14'd12171: ff_rdata <= 8'h00;
			14'd12172: ff_rdata <= 8'h45;
			14'd12173: ff_rdata <= 8'h6C;
			14'd12174: ff_rdata <= 8'h65;
			14'd12175: ff_rdata <= 8'h63;
			14'd12176: ff_rdata <= 8'h70;
			14'd12177: ff_rdata <= 8'h69;
			14'd12178: ff_rdata <= 8'h61;
			14'd12179: ff_rdata <= 8'h6E;
			14'd12180: ff_rdata <= 8'h00;
			14'd12181: ff_rdata <= 8'hED;
			14'd12182: ff_rdata <= 8'h0E;
			14'd12183: ff_rdata <= 8'h00;
			14'd12184: ff_rdata <= 8'h00;
			14'd12185: ff_rdata <= 8'h00;
			14'd12186: ff_rdata <= 8'h00;
			14'd12187: ff_rdata <= 8'h00;
			14'd12188: ff_rdata <= 8'h23;
			14'd12189: ff_rdata <= 8'h0F;
			14'd12190: ff_rdata <= 8'hDD;
			14'd12191: ff_rdata <= 8'h4A;
			14'd12192: ff_rdata <= 8'h20;
			14'd12193: ff_rdata <= 8'h00;
			14'd12194: ff_rdata <= 8'h00;
			14'd12195: ff_rdata <= 8'h00;
			14'd12196: ff_rdata <= 8'h43;
			14'd12197: ff_rdata <= 8'h00;
			14'd12198: ff_rdata <= 8'hBF;
			14'd12199: ff_rdata <= 8'h05;
			14'd12200: ff_rdata <= 8'h50;
			14'd12201: ff_rdata <= 8'h00;
			14'd12202: ff_rdata <= 8'h00;
			14'd12203: ff_rdata <= 8'h00;
			14'd12204: ff_rdata <= 8'h43;
			14'd12205: ff_rdata <= 8'h6C;
			14'd12206: ff_rdata <= 8'h61;
			14'd12207: ff_rdata <= 8'h76;
			14'd12208: ff_rdata <= 8'h69;
			14'd12209: ff_rdata <= 8'h63;
			14'd12210: ff_rdata <= 8'h6F;
			14'd12211: ff_rdata <= 8'h64;
			14'd12212: ff_rdata <= 8'h00;
			14'd12213: ff_rdata <= 8'hED;
			14'd12214: ff_rdata <= 8'h0C;
			14'd12215: ff_rdata <= 8'h00;
			14'd12216: ff_rdata <= 8'h00;
			14'd12217: ff_rdata <= 8'h00;
			14'd12218: ff_rdata <= 8'h00;
			14'd12219: ff_rdata <= 8'h00;
			14'd12220: ff_rdata <= 8'h03;
			14'd12221: ff_rdata <= 8'h11;
			14'd12222: ff_rdata <= 8'hD2;
			14'd12223: ff_rdata <= 8'hF4;
			14'd12224: ff_rdata <= 8'h20;
			14'd12225: ff_rdata <= 8'h00;
			14'd12226: ff_rdata <= 8'h00;
			14'd12227: ff_rdata <= 8'h00;
			14'd12228: ff_rdata <= 8'h09;
			14'd12229: ff_rdata <= 8'h08;
			14'd12230: ff_rdata <= 8'hB4;
			14'd12231: ff_rdata <= 8'hF5;
			14'd12232: ff_rdata <= 8'h60;
			14'd12233: ff_rdata <= 8'h00;
			14'd12234: ff_rdata <= 8'h00;
			14'd12235: ff_rdata <= 8'h00;
			14'd12236: ff_rdata <= 8'h48;
			14'd12237: ff_rdata <= 8'h61;
			14'd12238: ff_rdata <= 8'h72;
			14'd12239: ff_rdata <= 8'h70;
			14'd12240: ff_rdata <= 8'h73;
			14'd12241: ff_rdata <= 8'h69;
			14'd12242: ff_rdata <= 8'h63;
			14'd12243: ff_rdata <= 8'h64;
			14'd12244: ff_rdata <= 8'h00;
			14'd12245: ff_rdata <= 8'h0C;
			14'd12246: ff_rdata <= 8'h0D;
			14'd12247: ff_rdata <= 8'h00;
			14'd12248: ff_rdata <= 8'h00;
			14'd12249: ff_rdata <= 8'h00;
			14'd12250: ff_rdata <= 8'h00;
			14'd12251: ff_rdata <= 8'h00;
			14'd12252: ff_rdata <= 8'h01;
			14'd12253: ff_rdata <= 8'h06;
			14'd12254: ff_rdata <= 8'hA3;
			14'd12255: ff_rdata <= 8'hF4;
			14'd12256: ff_rdata <= 8'h40;
			14'd12257: ff_rdata <= 8'h00;
			14'd12258: ff_rdata <= 8'h00;
			14'd12259: ff_rdata <= 8'h00;
			14'd12260: ff_rdata <= 8'h00;
			14'd12261: ff_rdata <= 8'h19;
			14'd12262: ff_rdata <= 8'hE2;
			14'd12263: ff_rdata <= 8'hF4;
			14'd12264: ff_rdata <= 8'h00;
			14'd12265: ff_rdata <= 8'h00;
			14'd12266: ff_rdata <= 8'h00;
			14'd12267: ff_rdata <= 8'h00;
			14'd12268: ff_rdata <= 8'h48;
			14'd12269: ff_rdata <= 8'h61;
			14'd12270: ff_rdata <= 8'h72;
			14'd12271: ff_rdata <= 8'h70;
			14'd12272: ff_rdata <= 8'h73;
			14'd12273: ff_rdata <= 8'h63;
			14'd12274: ff_rdata <= 8'h64;
			14'd12275: ff_rdata <= 8'h32;
			14'd12276: ff_rdata <= 8'h00;
			14'd12277: ff_rdata <= 8'h00;
			14'd12278: ff_rdata <= 8'h0C;
			14'd12279: ff_rdata <= 8'h00;
			14'd12280: ff_rdata <= 8'h00;
			14'd12281: ff_rdata <= 8'h00;
			14'd12282: ff_rdata <= 8'h00;
			14'd12283: ff_rdata <= 8'h00;
			14'd12284: ff_rdata <= 8'h01;
			14'd12285: ff_rdata <= 8'h11;
			14'd12286: ff_rdata <= 8'hC0;
			14'd12287: ff_rdata <= 8'h01;
			14'd12288: ff_rdata <= 8'h20;
			14'd12289: ff_rdata <= 8'h00;
			14'd12290: ff_rdata <= 8'h00;
			14'd12291: ff_rdata <= 8'h00;
			14'd12292: ff_rdata <= 8'h01;
			14'd12293: ff_rdata <= 8'h08;
			14'd12294: ff_rdata <= 8'hB4;
			14'd12295: ff_rdata <= 8'hF6;
			14'd12296: ff_rdata <= 8'h80;
			14'd12297: ff_rdata <= 8'h00;
			14'd12298: ff_rdata <= 8'h00;
			14'd12299: ff_rdata <= 8'h00;
			14'd12300: ff_rdata <= 8'h56;
			14'd12301: ff_rdata <= 8'h69;
			14'd12302: ff_rdata <= 8'h62;
			14'd12303: ff_rdata <= 8'h72;
			14'd12304: ff_rdata <= 8'h61;
			14'd12305: ff_rdata <= 8'h70;
			14'd12306: ff_rdata <= 8'h68;
			14'd12307: ff_rdata <= 8'h6E;
			14'd12308: ff_rdata <= 8'h00;
			14'd12309: ff_rdata <= 8'h00;
			14'd12310: ff_rdata <= 8'hEC;
			14'd12311: ff_rdata <= 8'h00;
			14'd12312: ff_rdata <= 8'h00;
			14'd12313: ff_rdata <= 8'h00;
			14'd12314: ff_rdata <= 8'h00;
			14'd12315: ff_rdata <= 8'h00;
			14'd12316: ff_rdata <= 8'hF9;
			14'd12317: ff_rdata <= 8'h24;
			14'd12318: ff_rdata <= 8'h95;
			14'd12319: ff_rdata <= 8'hE5;
			14'd12320: ff_rdata <= 8'h80;
			14'd12321: ff_rdata <= 8'h00;
			14'd12322: ff_rdata <= 8'h00;
			14'd12323: ff_rdata <= 8'h00;
			14'd12324: ff_rdata <= 8'hF1;
			14'd12325: ff_rdata <= 8'h00;
			14'd12326: ff_rdata <= 8'hD1;
			14'd12327: ff_rdata <= 8'hF2;
			14'd12328: ff_rdata <= 8'h70;
			14'd12329: ff_rdata <= 8'h00;
			14'd12330: ff_rdata <= 8'h00;
			14'd12331: ff_rdata <= 8'h00;
			14'd12332: ff_rdata <= 8'h4B;
			14'd12333: ff_rdata <= 8'h6F;
			14'd12334: ff_rdata <= 8'h74;
			14'd12335: ff_rdata <= 8'h6F;
			14'd12336: ff_rdata <= 8'h20;
			14'd12337: ff_rdata <= 8'h20;
			14'd12338: ff_rdata <= 8'h20;
			14'd12339: ff_rdata <= 8'h20;
			14'd12340: ff_rdata <= 8'h00;
			14'd12341: ff_rdata <= 8'h00;
			14'd12342: ff_rdata <= 8'h0C;
			14'd12343: ff_rdata <= 8'h00;
			14'd12344: ff_rdata <= 8'h00;
			14'd12345: ff_rdata <= 8'h00;
			14'd12346: ff_rdata <= 8'h00;
			14'd12347: ff_rdata <= 8'h00;
			14'd12348: ff_rdata <= 8'h13;
			14'd12349: ff_rdata <= 8'h0C;
			14'd12350: ff_rdata <= 8'hFC;
			14'd12351: ff_rdata <= 8'h33;
			14'd12352: ff_rdata <= 8'h30;
			14'd12353: ff_rdata <= 8'h00;
			14'd12354: ff_rdata <= 8'h00;
			14'd12355: ff_rdata <= 8'h00;
			14'd12356: ff_rdata <= 8'h11;
			14'd12357: ff_rdata <= 8'h00;
			14'd12358: ff_rdata <= 8'hD2;
			14'd12359: ff_rdata <= 8'h83;
			14'd12360: ff_rdata <= 8'h80;
			14'd12361: ff_rdata <= 8'h00;
			14'd12362: ff_rdata <= 8'h00;
			14'd12363: ff_rdata <= 8'h00;
			14'd12364: ff_rdata <= 8'h54;
			14'd12365: ff_rdata <= 8'h61;
			14'd12366: ff_rdata <= 8'h69;
			14'd12367: ff_rdata <= 8'h6B;
			14'd12368: ff_rdata <= 8'h6F;
			14'd12369: ff_rdata <= 8'h20;
			14'd12370: ff_rdata <= 8'h20;
			14'd12371: ff_rdata <= 8'h20;
			14'd12372: ff_rdata <= 8'h00;
			14'd12373: ff_rdata <= 8'hF4;
			14'd12374: ff_rdata <= 8'h0E;
			14'd12375: ff_rdata <= 8'h00;
			14'd12376: ff_rdata <= 8'h00;
			14'd12377: ff_rdata <= 8'h00;
			14'd12378: ff_rdata <= 8'h00;
			14'd12379: ff_rdata <= 8'h00;
			14'd12380: ff_rdata <= 8'h01;
			14'd12381: ff_rdata <= 8'h0E;
			14'd12382: ff_rdata <= 8'hCA;
			14'd12383: ff_rdata <= 8'h44;
			14'd12384: ff_rdata <= 8'h20;
			14'd12385: ff_rdata <= 8'h00;
			14'd12386: ff_rdata <= 8'h00;
			14'd12387: ff_rdata <= 8'h00;
			14'd12388: ff_rdata <= 8'h10;
			14'd12389: ff_rdata <= 8'h00;
			14'd12390: ff_rdata <= 8'hE6;
			14'd12391: ff_rdata <= 8'h24;
			14'd12392: ff_rdata <= 8'h80;
			14'd12393: ff_rdata <= 8'h00;
			14'd12394: ff_rdata <= 8'h00;
			14'd12395: ff_rdata <= 8'h00;
			14'd12396: ff_rdata <= 8'h45;
			14'd12397: ff_rdata <= 8'h6E;
			14'd12398: ff_rdata <= 8'h67;
			14'd12399: ff_rdata <= 8'h69;
			14'd12400: ff_rdata <= 8'h6E;
			14'd12401: ff_rdata <= 8'h65;
			14'd12402: ff_rdata <= 8'h20;
			14'd12403: ff_rdata <= 8'h20;
			14'd12404: ff_rdata <= 8'h00;
			14'd12405: ff_rdata <= 8'hE8;
			14'd12406: ff_rdata <= 8'h6E;
			14'd12407: ff_rdata <= 8'h00;
			14'd12408: ff_rdata <= 8'h00;
			14'd12409: ff_rdata <= 8'h00;
			14'd12410: ff_rdata <= 8'h00;
			14'd12411: ff_rdata <= 8'h00;
			14'd12412: ff_rdata <= 8'hE0;
			14'd12413: ff_rdata <= 8'h1B;
			14'd12414: ff_rdata <= 8'h11;
			14'd12415: ff_rdata <= 8'h04;
			14'd12416: ff_rdata <= 8'h40;
			14'd12417: ff_rdata <= 8'h00;
			14'd12418: ff_rdata <= 8'h00;
			14'd12419: ff_rdata <= 8'h00;
			14'd12420: ff_rdata <= 8'hF4;
			14'd12421: ff_rdata <= 8'h80;
			14'd12422: ff_rdata <= 8'hF0;
			14'd12423: ff_rdata <= 8'h08;
			14'd12424: ff_rdata <= 8'h50;
			14'd12425: ff_rdata <= 8'h00;
			14'd12426: ff_rdata <= 8'h00;
			14'd12427: ff_rdata <= 8'h00;
			14'd12428: ff_rdata <= 8'h55;
			14'd12429: ff_rdata <= 8'h46;
			14'd12430: ff_rdata <= 8'h4F;
			14'd12431: ff_rdata <= 8'h20;
			14'd12432: ff_rdata <= 8'h20;
			14'd12433: ff_rdata <= 8'h20;
			14'd12434: ff_rdata <= 8'h20;
			14'd12435: ff_rdata <= 8'h20;
			14'd12436: ff_rdata <= 8'h00;
			14'd12437: ff_rdata <= 8'h0C;
			14'd12438: ff_rdata <= 8'hEE;
			14'd12439: ff_rdata <= 8'h00;
			14'd12440: ff_rdata <= 8'h00;
			14'd12441: ff_rdata <= 8'h00;
			14'd12442: ff_rdata <= 8'h00;
			14'd12443: ff_rdata <= 8'h00;
			14'd12444: ff_rdata <= 8'hFF;
			14'd12445: ff_rdata <= 8'h19;
			14'd12446: ff_rdata <= 8'h50;
			14'd12447: ff_rdata <= 8'h05;
			14'd12448: ff_rdata <= 8'h60;
			14'd12449: ff_rdata <= 8'h00;
			14'd12450: ff_rdata <= 8'h00;
			14'd12451: ff_rdata <= 8'h00;
			14'd12452: ff_rdata <= 8'h70;
			14'd12453: ff_rdata <= 8'h00;
			14'd12454: ff_rdata <= 8'h1F;
			14'd12455: ff_rdata <= 8'h01;
			14'd12456: ff_rdata <= 8'h40;
			14'd12457: ff_rdata <= 8'h00;
			14'd12458: ff_rdata <= 8'h00;
			14'd12459: ff_rdata <= 8'h00;
			14'd12460: ff_rdata <= 8'h53;
			14'd12461: ff_rdata <= 8'h79;
			14'd12462: ff_rdata <= 8'h6E;
			14'd12463: ff_rdata <= 8'h42;
			14'd12464: ff_rdata <= 8'h65;
			14'd12465: ff_rdata <= 8'h6C;
			14'd12466: ff_rdata <= 8'h6C;
			14'd12467: ff_rdata <= 8'h20;
			14'd12468: ff_rdata <= 8'h00;
			14'd12469: ff_rdata <= 8'h00;
			14'd12470: ff_rdata <= 8'h0E;
			14'd12471: ff_rdata <= 8'h00;
			14'd12472: ff_rdata <= 8'h00;
			14'd12473: ff_rdata <= 8'h00;
			14'd12474: ff_rdata <= 8'h00;
			14'd12475: ff_rdata <= 8'h00;
			14'd12476: ff_rdata <= 8'h13;
			14'd12477: ff_rdata <= 8'h11;
			14'd12478: ff_rdata <= 8'hFA;
			14'd12479: ff_rdata <= 8'h21;
			14'd12480: ff_rdata <= 8'h30;
			14'd12481: ff_rdata <= 8'h00;
			14'd12482: ff_rdata <= 8'h00;
			14'd12483: ff_rdata <= 8'h00;
			14'd12484: ff_rdata <= 8'h11;
			14'd12485: ff_rdata <= 8'h00;
			14'd12486: ff_rdata <= 8'hF2;
			14'd12487: ff_rdata <= 8'hF4;
			14'd12488: ff_rdata <= 8'h80;
			14'd12489: ff_rdata <= 8'h00;
			14'd12490: ff_rdata <= 8'h00;
			14'd12491: ff_rdata <= 8'h00;
			14'd12492: ff_rdata <= 8'h43;
			14'd12493: ff_rdata <= 8'h68;
			14'd12494: ff_rdata <= 8'h69;
			14'd12495: ff_rdata <= 8'h6D;
			14'd12496: ff_rdata <= 8'h65;
			14'd12497: ff_rdata <= 8'h20;
			14'd12498: ff_rdata <= 8'h20;
			14'd12499: ff_rdata <= 8'h20;
			14'd12500: ff_rdata <= 8'h00;
			14'd12501: ff_rdata <= 8'h00;
			14'd12502: ff_rdata <= 8'hEA;
			14'd12503: ff_rdata <= 8'h00;
			14'd12504: ff_rdata <= 8'h00;
			14'd12505: ff_rdata <= 8'h00;
			14'd12506: ff_rdata <= 8'h00;
			14'd12507: ff_rdata <= 8'h00;
			14'd12508: ff_rdata <= 8'hA6;
			14'd12509: ff_rdata <= 8'h10;
			14'd12510: ff_rdata <= 8'hFB;
			14'd12511: ff_rdata <= 8'h11;
			14'd12512: ff_rdata <= 8'h20;
			14'd12513: ff_rdata <= 8'h00;
			14'd12514: ff_rdata <= 8'h00;
			14'd12515: ff_rdata <= 8'h00;
			14'd12516: ff_rdata <= 8'h42;
			14'd12517: ff_rdata <= 8'h0B;
			14'd12518: ff_rdata <= 8'hB9;
			14'd12519: ff_rdata <= 8'h02;
			14'd12520: ff_rdata <= 8'h60;
			14'd12521: ff_rdata <= 8'h00;
			14'd12522: ff_rdata <= 8'h00;
			14'd12523: ff_rdata <= 8'h00;
			14'd12524: ff_rdata <= 8'h53;
			14'd12525: ff_rdata <= 8'h79;
			14'd12526: ff_rdata <= 8'h6E;
			14'd12527: ff_rdata <= 8'h42;
			14'd12528: ff_rdata <= 8'h61;
			14'd12529: ff_rdata <= 8'h73;
			14'd12530: ff_rdata <= 8'h73;
			14'd12531: ff_rdata <= 8'h20;
			14'd12532: ff_rdata <= 8'hF8;
			14'd12533: ff_rdata <= 8'hF3;
			14'd12534: ff_rdata <= 8'h0C;
			14'd12535: ff_rdata <= 8'h00;
			14'd12536: ff_rdata <= 8'h00;
			14'd12537: ff_rdata <= 8'h00;
			14'd12538: ff_rdata <= 8'h00;
			14'd12539: ff_rdata <= 8'h00;
			14'd12540: ff_rdata <= 8'h40;
			14'd12541: ff_rdata <= 8'h89;
			14'd12542: ff_rdata <= 8'hC7;
			14'd12543: ff_rdata <= 8'h14;
			14'd12544: ff_rdata <= 8'h40;
			14'd12545: ff_rdata <= 8'h00;
			14'd12546: ff_rdata <= 8'h00;
			14'd12547: ff_rdata <= 8'h00;
			14'd12548: ff_rdata <= 8'h31;
			14'd12549: ff_rdata <= 8'h00;
			14'd12550: ff_rdata <= 8'hF9;
			14'd12551: ff_rdata <= 8'h04;
			14'd12552: ff_rdata <= 8'h80;
			14'd12553: ff_rdata <= 8'h00;
			14'd12554: ff_rdata <= 8'h00;
			14'd12555: ff_rdata <= 8'h00;
			14'd12556: ff_rdata <= 8'h53;
			14'd12557: ff_rdata <= 8'h79;
			14'd12558: ff_rdata <= 8'h6E;
			14'd12559: ff_rdata <= 8'h74;
			14'd12560: ff_rdata <= 8'h68;
			14'd12561: ff_rdata <= 8'h73;
			14'd12562: ff_rdata <= 8'h69;
			14'd12563: ff_rdata <= 8'h7A;
			14'd12564: ff_rdata <= 8'h00;
			14'd12565: ff_rdata <= 8'hE8;
			14'd12566: ff_rdata <= 8'h6C;
			14'd12567: ff_rdata <= 8'h00;
			14'd12568: ff_rdata <= 8'h00;
			14'd12569: ff_rdata <= 8'h00;
			14'd12570: ff_rdata <= 8'h00;
			14'd12571: ff_rdata <= 8'h00;
			14'd12572: ff_rdata <= 8'h42;
			14'd12573: ff_rdata <= 8'h0B;
			14'd12574: ff_rdata <= 8'h94;
			14'd12575: ff_rdata <= 8'h33;
			14'd12576: ff_rdata <= 8'h00;
			14'd12577: ff_rdata <= 8'h00;
			14'd12578: ff_rdata <= 8'h00;
			14'd12579: ff_rdata <= 8'h00;
			14'd12580: ff_rdata <= 8'h44;
			14'd12581: ff_rdata <= 8'h05;
			14'd12582: ff_rdata <= 8'hB0;
			14'd12583: ff_rdata <= 8'hF6;
			14'd12584: ff_rdata <= 8'h50;
			14'd12585: ff_rdata <= 8'h00;
			14'd12586: ff_rdata <= 8'h00;
			14'd12587: ff_rdata <= 8'h00;
			14'd12588: ff_rdata <= 8'h53;
			14'd12589: ff_rdata <= 8'h79;
			14'd12590: ff_rdata <= 8'h6E;
			14'd12591: ff_rdata <= 8'h50;
			14'd12592: ff_rdata <= 8'h65;
			14'd12593: ff_rdata <= 8'h72;
			14'd12594: ff_rdata <= 8'h63;
			14'd12595: ff_rdata <= 8'h75;
			14'd12596: ff_rdata <= 8'h00;
			14'd12597: ff_rdata <= 8'hF4;
			14'd12598: ff_rdata <= 8'h0E;
			14'd12599: ff_rdata <= 8'h00;
			14'd12600: ff_rdata <= 8'h00;
			14'd12601: ff_rdata <= 8'h00;
			14'd12602: ff_rdata <= 8'h00;
			14'd12603: ff_rdata <= 8'h00;
			14'd12604: ff_rdata <= 8'h01;
			14'd12605: ff_rdata <= 8'h0B;
			14'd12606: ff_rdata <= 8'hBA;
			14'd12607: ff_rdata <= 8'h25;
			14'd12608: ff_rdata <= 8'h60;
			14'd12609: ff_rdata <= 8'h00;
			14'd12610: ff_rdata <= 8'h00;
			14'd12611: ff_rdata <= 8'h00;
			14'd12612: ff_rdata <= 8'h03;
			14'd12613: ff_rdata <= 8'h00;
			14'd12614: ff_rdata <= 8'hD9;
			14'd12615: ff_rdata <= 8'h06;
			14'd12616: ff_rdata <= 8'h80;
			14'd12617: ff_rdata <= 8'h00;
			14'd12618: ff_rdata <= 8'h00;
			14'd12619: ff_rdata <= 8'h00;
			14'd12620: ff_rdata <= 8'h53;
			14'd12621: ff_rdata <= 8'h79;
			14'd12622: ff_rdata <= 8'h6E;
			14'd12623: ff_rdata <= 8'h52;
			14'd12624: ff_rdata <= 8'h68;
			14'd12625: ff_rdata <= 8'h79;
			14'd12626: ff_rdata <= 8'h74;
			14'd12627: ff_rdata <= 8'h68;
			14'd12628: ff_rdata <= 8'h00;
			14'd12629: ff_rdata <= 8'h0C;
			14'd12630: ff_rdata <= 8'h0E;
			14'd12631: ff_rdata <= 8'h00;
			14'd12632: ff_rdata <= 8'h00;
			14'd12633: ff_rdata <= 8'h00;
			14'd12634: ff_rdata <= 8'h00;
			14'd12635: ff_rdata <= 8'h00;
			14'd12636: ff_rdata <= 8'h40;
			14'd12637: ff_rdata <= 8'h00;
			14'd12638: ff_rdata <= 8'hFA;
			14'd12639: ff_rdata <= 8'h37;
			14'd12640: ff_rdata <= 8'h40;
			14'd12641: ff_rdata <= 8'h00;
			14'd12642: ff_rdata <= 8'h00;
			14'd12643: ff_rdata <= 8'h00;
			14'd12644: ff_rdata <= 8'h00;
			14'd12645: ff_rdata <= 8'h00;
			14'd12646: ff_rdata <= 8'hD9;
			14'd12647: ff_rdata <= 8'h04;
			14'd12648: ff_rdata <= 8'h00;
			14'd12649: ff_rdata <= 8'h00;
			14'd12650: ff_rdata <= 8'h00;
			14'd12651: ff_rdata <= 8'h00;
			14'd12652: ff_rdata <= 8'h48;
			14'd12653: ff_rdata <= 8'h61;
			14'd12654: ff_rdata <= 8'h72;
			14'd12655: ff_rdata <= 8'h6D;
			14'd12656: ff_rdata <= 8'h44;
			14'd12657: ff_rdata <= 8'h72;
			14'd12658: ff_rdata <= 8'h75;
			14'd12659: ff_rdata <= 8'h6D;
			14'd12660: ff_rdata <= 8'h00;
			14'd12661: ff_rdata <= 8'hE1;
			14'd12662: ff_rdata <= 8'h0E;
			14'd12663: ff_rdata <= 8'h00;
			14'd12664: ff_rdata <= 8'h00;
			14'd12665: ff_rdata <= 8'h00;
			14'd12666: ff_rdata <= 8'h00;
			14'd12667: ff_rdata <= 8'h00;
			14'd12668: ff_rdata <= 8'h02;
			14'd12669: ff_rdata <= 8'h09;
			14'd12670: ff_rdata <= 8'hCB;
			14'd12671: ff_rdata <= 8'h39;
			14'd12672: ff_rdata <= 8'h60;
			14'd12673: ff_rdata <= 8'h00;
			14'd12674: ff_rdata <= 8'h00;
			14'd12675: ff_rdata <= 8'h00;
			14'd12676: ff_rdata <= 8'h03;
			14'd12677: ff_rdata <= 8'h00;
			14'd12678: ff_rdata <= 8'hFF;
			14'd12679: ff_rdata <= 8'h06;
			14'd12680: ff_rdata <= 8'h80;
			14'd12681: ff_rdata <= 8'h00;
			14'd12682: ff_rdata <= 8'h00;
			14'd12683: ff_rdata <= 8'h00;
			14'd12684: ff_rdata <= 8'h43;
			14'd12685: ff_rdata <= 8'h6F;
			14'd12686: ff_rdata <= 8'h77;
			14'd12687: ff_rdata <= 8'h62;
			14'd12688: ff_rdata <= 8'h65;
			14'd12689: ff_rdata <= 8'h6C;
			14'd12690: ff_rdata <= 8'h6C;
			14'd12691: ff_rdata <= 8'h20;
			14'd12692: ff_rdata <= 8'h00;
			14'd12693: ff_rdata <= 8'hF4;
			14'd12694: ff_rdata <= 8'h0A;
			14'd12695: ff_rdata <= 8'h00;
			14'd12696: ff_rdata <= 8'h00;
			14'd12697: ff_rdata <= 8'h00;
			14'd12698: ff_rdata <= 8'h00;
			14'd12699: ff_rdata <= 8'h00;
			14'd12700: ff_rdata <= 8'h18;
			14'd12701: ff_rdata <= 8'h09;
			14'd12702: ff_rdata <= 8'hF8;
			14'd12703: ff_rdata <= 8'h26;
			14'd12704: ff_rdata <= 8'h20;
			14'd12705: ff_rdata <= 8'h00;
			14'd12706: ff_rdata <= 8'h00;
			14'd12707: ff_rdata <= 8'h00;
			14'd12708: ff_rdata <= 8'h11;
			14'd12709: ff_rdata <= 8'h00;
			14'd12710: ff_rdata <= 8'hF5;
			14'd12711: ff_rdata <= 8'h26;
			14'd12712: ff_rdata <= 8'h60;
			14'd12713: ff_rdata <= 8'h00;
			14'd12714: ff_rdata <= 8'h00;
			14'd12715: ff_rdata <= 8'h00;
			14'd12716: ff_rdata <= 8'h43;
			14'd12717: ff_rdata <= 8'h6C;
			14'd12718: ff_rdata <= 8'h73;
			14'd12719: ff_rdata <= 8'h65;
			14'd12720: ff_rdata <= 8'h48;
			14'd12721: ff_rdata <= 8'h69;
			14'd12722: ff_rdata <= 8'h68;
			14'd12723: ff_rdata <= 8'h74;
			14'd12724: ff_rdata <= 8'h00;
			14'd12725: ff_rdata <= 8'h18;
			14'd12726: ff_rdata <= 8'h0E;
			14'd12727: ff_rdata <= 8'h00;
			14'd12728: ff_rdata <= 8'h00;
			14'd12729: ff_rdata <= 8'h00;
			14'd12730: ff_rdata <= 8'h00;
			14'd12731: ff_rdata <= 8'h00;
			14'd12732: ff_rdata <= 8'h0B;
			14'd12733: ff_rdata <= 8'h09;
			14'd12734: ff_rdata <= 8'hF0;
			14'd12735: ff_rdata <= 8'h01;
			14'd12736: ff_rdata <= 8'h80;
			14'd12737: ff_rdata <= 8'h00;
			14'd12738: ff_rdata <= 8'h00;
			14'd12739: ff_rdata <= 8'h00;
			14'd12740: ff_rdata <= 8'h04;
			14'd12741: ff_rdata <= 8'h00;
			14'd12742: ff_rdata <= 8'hF5;
			14'd12743: ff_rdata <= 8'h27;
			14'd12744: ff_rdata <= 8'h80;
			14'd12745: ff_rdata <= 8'h00;
			14'd12746: ff_rdata <= 8'h00;
			14'd12747: ff_rdata <= 8'h00;
			14'd12748: ff_rdata <= 8'h53;
			14'd12749: ff_rdata <= 8'h6E;
			14'd12750: ff_rdata <= 8'h61;
			14'd12751: ff_rdata <= 8'h72;
			14'd12752: ff_rdata <= 8'h65;
			14'd12753: ff_rdata <= 8'h44;
			14'd12754: ff_rdata <= 8'h72;
			14'd12755: ff_rdata <= 8'h6D;
			14'd12756: ff_rdata <= 8'h00;
			14'd12757: ff_rdata <= 8'h00;
			14'd12758: ff_rdata <= 8'h6E;
			14'd12759: ff_rdata <= 8'h00;
			14'd12760: ff_rdata <= 8'h00;
			14'd12761: ff_rdata <= 8'h00;
			14'd12762: ff_rdata <= 8'h00;
			14'd12763: ff_rdata <= 8'h00;
			14'd12764: ff_rdata <= 8'h40;
			14'd12765: ff_rdata <= 8'h07;
			14'd12766: ff_rdata <= 8'hD0;
			14'd12767: ff_rdata <= 8'h01;
			14'd12768: ff_rdata <= 8'h80;
			14'd12769: ff_rdata <= 8'h00;
			14'd12770: ff_rdata <= 8'h00;
			14'd12771: ff_rdata <= 8'h00;
			14'd12772: ff_rdata <= 8'h40;
			14'd12773: ff_rdata <= 8'h00;
			14'd12774: ff_rdata <= 8'hD6;
			14'd12775: ff_rdata <= 8'h27;
			14'd12776: ff_rdata <= 8'h80;
			14'd12777: ff_rdata <= 8'h00;
			14'd12778: ff_rdata <= 8'h00;
			14'd12779: ff_rdata <= 8'h00;
			14'd12780: ff_rdata <= 8'h42;
			14'd12781: ff_rdata <= 8'h61;
			14'd12782: ff_rdata <= 8'h73;
			14'd12783: ff_rdata <= 8'h73;
			14'd12784: ff_rdata <= 8'h44;
			14'd12785: ff_rdata <= 8'h72;
			14'd12786: ff_rdata <= 8'h75;
			14'd12787: ff_rdata <= 8'h6D;
			14'd12788: ff_rdata <= 8'h00;
			14'd12789: ff_rdata <= 8'hF4;
			14'd12790: ff_rdata <= 8'h0C;
			14'd12791: ff_rdata <= 8'h00;
			14'd12792: ff_rdata <= 8'h00;
			14'd12793: ff_rdata <= 8'h00;
			14'd12794: ff_rdata <= 8'h00;
			14'd12795: ff_rdata <= 8'h00;
			14'd12796: ff_rdata <= 8'h00;
			14'd12797: ff_rdata <= 8'h07;
			14'd12798: ff_rdata <= 8'hCB;
			14'd12799: ff_rdata <= 8'h36;
			14'd12800: ff_rdata <= 8'h40;
			14'd12801: ff_rdata <= 8'h00;
			14'd12802: ff_rdata <= 8'h00;
			14'd12803: ff_rdata <= 8'h00;
			14'd12804: ff_rdata <= 8'h01;
			14'd12805: ff_rdata <= 8'h00;
			14'd12806: ff_rdata <= 8'hE3;
			14'd12807: ff_rdata <= 8'h25;
			14'd12808: ff_rdata <= 8'h80;
			14'd12809: ff_rdata <= 8'h00;
			14'd12810: ff_rdata <= 8'h00;
			14'd12811: ff_rdata <= 8'h00;
			14'd12812: ff_rdata <= 8'h50;
			14'd12813: ff_rdata <= 8'h69;
			14'd12814: ff_rdata <= 8'h61;
			14'd12815: ff_rdata <= 8'h6E;
			14'd12816: ff_rdata <= 8'h6F;
			14'd12817: ff_rdata <= 8'h20;
			14'd12818: ff_rdata <= 8'h33;
			14'd12819: ff_rdata <= 8'h20;
			14'd12820: ff_rdata <= 8'h00;
			14'd12821: ff_rdata <= 8'h00;
			14'd12822: ff_rdata <= 8'h08;
			14'd12823: ff_rdata <= 8'h00;
			14'd12824: ff_rdata <= 8'h00;
			14'd12825: ff_rdata <= 8'h00;
			14'd12826: ff_rdata <= 8'h00;
			14'd12827: ff_rdata <= 8'h00;
			14'd12828: ff_rdata <= 8'h11;
			14'd12829: ff_rdata <= 8'h08;
			14'd12830: ff_rdata <= 8'hFA;
			14'd12831: ff_rdata <= 8'h20;
			14'd12832: ff_rdata <= 8'h30;
			14'd12833: ff_rdata <= 8'h00;
			14'd12834: ff_rdata <= 8'h00;
			14'd12835: ff_rdata <= 8'h00;
			14'd12836: ff_rdata <= 8'h11;
			14'd12837: ff_rdata <= 8'h00;
			14'd12838: ff_rdata <= 8'hB2;
			14'd12839: ff_rdata <= 8'hF4;
			14'd12840: ff_rdata <= 8'h70;
			14'd12841: ff_rdata <= 8'h00;
			14'd12842: ff_rdata <= 8'h00;
			14'd12843: ff_rdata <= 8'h00;
			14'd12844: ff_rdata <= 8'h45;
			14'd12845: ff_rdata <= 8'h6C;
			14'd12846: ff_rdata <= 8'h65;
			14'd12847: ff_rdata <= 8'h63;
			14'd12848: ff_rdata <= 8'h70;
			14'd12849: ff_rdata <= 8'h69;
			14'd12850: ff_rdata <= 8'h61;
			14'd12851: ff_rdata <= 8'h32;
			14'd12852: ff_rdata <= 8'h00;
			14'd12853: ff_rdata <= 8'h00;
			14'd12854: ff_rdata <= 8'h00;
			14'd12855: ff_rdata <= 8'h00;
			14'd12856: ff_rdata <= 8'h00;
			14'd12857: ff_rdata <= 8'h00;
			14'd12858: ff_rdata <= 8'h00;
			14'd12859: ff_rdata <= 8'h00;
			14'd12860: ff_rdata <= 8'h11;
			14'd12861: ff_rdata <= 8'h11;
			14'd12862: ff_rdata <= 8'hC0;
			14'd12863: ff_rdata <= 8'h01;
			14'd12864: ff_rdata <= 8'h10;
			14'd12865: ff_rdata <= 8'h00;
			14'd12866: ff_rdata <= 8'h00;
			14'd12867: ff_rdata <= 8'h00;
			14'd12868: ff_rdata <= 8'h11;
			14'd12869: ff_rdata <= 8'h00;
			14'd12870: ff_rdata <= 8'hB2;
			14'd12871: ff_rdata <= 8'hF4;
			14'd12872: ff_rdata <= 8'h80;
			14'd12873: ff_rdata <= 8'h00;
			14'd12874: ff_rdata <= 8'h00;
			14'd12875: ff_rdata <= 8'h00;
			14'd12876: ff_rdata <= 8'h53;
			14'd12877: ff_rdata <= 8'h61;
			14'd12878: ff_rdata <= 8'h6E;
			14'd12879: ff_rdata <= 8'h74;
			14'd12880: ff_rdata <= 8'h6F;
			14'd12881: ff_rdata <= 8'h6F;
			14'd12882: ff_rdata <= 8'h6C;
			14'd12883: ff_rdata <= 8'h32;
			14'd12884: ff_rdata <= 8'h00;
			14'd12885: ff_rdata <= 8'hED;
			14'd12886: ff_rdata <= 8'h0E;
			14'd12887: ff_rdata <= 8'h00;
			14'd12888: ff_rdata <= 8'h00;
			14'd12889: ff_rdata <= 8'h00;
			14'd12890: ff_rdata <= 8'h00;
			14'd12891: ff_rdata <= 8'h00;
			14'd12892: ff_rdata <= 8'h19;
			14'd12893: ff_rdata <= 8'h15;
			14'd12894: ff_rdata <= 8'hE7;
			14'd12895: ff_rdata <= 8'h21;
			14'd12896: ff_rdata <= 8'h80;
			14'd12897: ff_rdata <= 8'h00;
			14'd12898: ff_rdata <= 8'h00;
			14'd12899: ff_rdata <= 8'h00;
			14'd12900: ff_rdata <= 8'h53;
			14'd12901: ff_rdata <= 8'h03;
			14'd12902: ff_rdata <= 8'h95;
			14'd12903: ff_rdata <= 8'h03;
			14'd12904: ff_rdata <= 8'h60;
			14'd12905: ff_rdata <= 8'h00;
			14'd12906: ff_rdata <= 8'h00;
			14'd12907: ff_rdata <= 8'h00;
			14'd12908: ff_rdata <= 8'h42;
			14'd12909: ff_rdata <= 8'h72;
			14'd12910: ff_rdata <= 8'h61;
			14'd12911: ff_rdata <= 8'h73;
			14'd12912: ff_rdata <= 8'h73;
			14'd12913: ff_rdata <= 8'h20;
			14'd12914: ff_rdata <= 8'h20;
			14'd12915: ff_rdata <= 8'h20;
			14'd12916: ff_rdata <= 8'h00;
			14'd12917: ff_rdata <= 8'h00;
			14'd12918: ff_rdata <= 8'h6E;
			14'd12919: ff_rdata <= 8'h00;
			14'd12920: ff_rdata <= 8'h00;
			14'd12921: ff_rdata <= 8'h00;
			14'd12922: ff_rdata <= 8'h00;
			14'd12923: ff_rdata <= 8'h00;
			14'd12924: ff_rdata <= 8'h30;
			14'd12925: ff_rdata <= 8'h19;
			14'd12926: ff_rdata <= 8'h42;
			14'd12927: ff_rdata <= 8'h26;
			14'd12928: ff_rdata <= 8'h40;
			14'd12929: ff_rdata <= 8'h00;
			14'd12930: ff_rdata <= 8'h00;
			14'd12931: ff_rdata <= 8'h00;
			14'd12932: ff_rdata <= 8'h70;
			14'd12933: ff_rdata <= 8'h00;
			14'd12934: ff_rdata <= 8'h62;
			14'd12935: ff_rdata <= 8'h24;
			14'd12936: ff_rdata <= 8'h60;
			14'd12937: ff_rdata <= 8'h00;
			14'd12938: ff_rdata <= 8'h00;
			14'd12939: ff_rdata <= 8'h00;
			14'd12940: ff_rdata <= 8'h46;
			14'd12941: ff_rdata <= 8'h6C;
			14'd12942: ff_rdata <= 8'h75;
			14'd12943: ff_rdata <= 8'h74;
			14'd12944: ff_rdata <= 8'h65;
			14'd12945: ff_rdata <= 8'h20;
			14'd12946: ff_rdata <= 8'h32;
			14'd12947: ff_rdata <= 8'h20;
			14'd12948: ff_rdata <= 8'h00;
			14'd12949: ff_rdata <= 8'h0C;
			14'd12950: ff_rdata <= 8'h0E;
			14'd12951: ff_rdata <= 8'h00;
			14'd12952: ff_rdata <= 8'h00;
			14'd12953: ff_rdata <= 8'h00;
			14'd12954: ff_rdata <= 8'h00;
			14'd12955: ff_rdata <= 8'h00;
			14'd12956: ff_rdata <= 8'h62;
			14'd12957: ff_rdata <= 8'h25;
			14'd12958: ff_rdata <= 8'h64;
			14'd12959: ff_rdata <= 8'h12;
			14'd12960: ff_rdata <= 8'h40;
			14'd12961: ff_rdata <= 8'h00;
			14'd12962: ff_rdata <= 8'h00;
			14'd12963: ff_rdata <= 8'h00;
			14'd12964: ff_rdata <= 8'h71;
			14'd12965: ff_rdata <= 8'h03;
			14'd12966: ff_rdata <= 8'h43;
			14'd12967: ff_rdata <= 8'h26;
			14'd12968: ff_rdata <= 8'h80;
			14'd12969: ff_rdata <= 8'h00;
			14'd12970: ff_rdata <= 8'h00;
			14'd12971: ff_rdata <= 8'h00;
			14'd12972: ff_rdata <= 8'h43;
			14'd12973: ff_rdata <= 8'h6C;
			14'd12974: ff_rdata <= 8'h61;
			14'd12975: ff_rdata <= 8'h76;
			14'd12976: ff_rdata <= 8'h69;
			14'd12977: ff_rdata <= 8'h63;
			14'd12978: ff_rdata <= 8'h64;
			14'd12979: ff_rdata <= 8'h32;
			14'd12980: ff_rdata <= 8'h00;
			14'd12981: ff_rdata <= 8'h0C;
			14'd12982: ff_rdata <= 8'h0A;
			14'd12983: ff_rdata <= 8'h00;
			14'd12984: ff_rdata <= 8'h00;
			14'd12985: ff_rdata <= 8'h00;
			14'd12986: ff_rdata <= 8'h00;
			14'd12987: ff_rdata <= 8'h00;
			14'd12988: ff_rdata <= 8'h21;
			14'd12989: ff_rdata <= 8'h0B;
			14'd12990: ff_rdata <= 8'h90;
			14'd12991: ff_rdata <= 8'h02;
			14'd12992: ff_rdata <= 8'h50;
			14'd12993: ff_rdata <= 8'h00;
			14'd12994: ff_rdata <= 8'h00;
			14'd12995: ff_rdata <= 8'h00;
			14'd12996: ff_rdata <= 8'h03;
			14'd12997: ff_rdata <= 8'h03;
			14'd12998: ff_rdata <= 8'hD4;
			14'd12999: ff_rdata <= 8'hF5;
			14'd13000: ff_rdata <= 8'h60;
			14'd13001: ff_rdata <= 8'h00;
			14'd13002: ff_rdata <= 8'h00;
			14'd13003: ff_rdata <= 8'h00;
			14'd13004: ff_rdata <= 8'h43;
			14'd13005: ff_rdata <= 8'h6C;
			14'd13006: ff_rdata <= 8'h61;
			14'd13007: ff_rdata <= 8'h76;
			14'd13008: ff_rdata <= 8'h69;
			14'd13009: ff_rdata <= 8'h63;
			14'd13010: ff_rdata <= 8'h64;
			14'd13011: ff_rdata <= 8'h33;
			14'd13012: ff_rdata <= 8'h00;
			14'd13013: ff_rdata <= 8'h0C;
			14'd13014: ff_rdata <= 8'h0A;
			14'd13015: ff_rdata <= 8'h00;
			14'd13016: ff_rdata <= 8'h00;
			14'd13017: ff_rdata <= 8'h00;
			14'd13018: ff_rdata <= 8'h00;
			14'd13019: ff_rdata <= 8'h00;
			14'd13020: ff_rdata <= 8'h01;
			14'd13021: ff_rdata <= 8'h0A;
			14'd13022: ff_rdata <= 8'h90;
			14'd13023: ff_rdata <= 8'h03;
			14'd13024: ff_rdata <= 8'h40;
			14'd13025: ff_rdata <= 8'h00;
			14'd13026: ff_rdata <= 8'h00;
			14'd13027: ff_rdata <= 8'h00;
			14'd13028: ff_rdata <= 8'h03;
			14'd13029: ff_rdata <= 8'h03;
			14'd13030: ff_rdata <= 8'hA4;
			14'd13031: ff_rdata <= 8'hF5;
			14'd13032: ff_rdata <= 8'h60;
			14'd13033: ff_rdata <= 8'h00;
			14'd13034: ff_rdata <= 8'h00;
			14'd13035: ff_rdata <= 8'h00;
			14'd13036: ff_rdata <= 8'h4B;
			14'd13037: ff_rdata <= 8'h6F;
			14'd13038: ff_rdata <= 8'h74;
			14'd13039: ff_rdata <= 8'h6F;
			14'd13040: ff_rdata <= 8'h20;
			14'd13041: ff_rdata <= 8'h32;
			14'd13042: ff_rdata <= 8'h20;
			14'd13043: ff_rdata <= 8'h20;
			14'd13044: ff_rdata <= 8'h00;
			14'd13045: ff_rdata <= 8'hED;
			14'd13046: ff_rdata <= 8'h0A;
			14'd13047: ff_rdata <= 8'h00;
			14'd13048: ff_rdata <= 8'h00;
			14'd13049: ff_rdata <= 8'h00;
			14'd13050: ff_rdata <= 8'h00;
			14'd13051: ff_rdata <= 8'h00;
			14'd13052: ff_rdata <= 8'h43;
			14'd13053: ff_rdata <= 8'h0E;
			14'd13054: ff_rdata <= 8'hB5;
			14'd13055: ff_rdata <= 8'h84;
			14'd13056: ff_rdata <= 8'h50;
			14'd13057: ff_rdata <= 8'h00;
			14'd13058: ff_rdata <= 8'h00;
			14'd13059: ff_rdata <= 8'h00;
			14'd13060: ff_rdata <= 8'h53;
			14'd13061: ff_rdata <= 8'h81;
			14'd13062: ff_rdata <= 8'hE9;
			14'd13063: ff_rdata <= 8'h04;
			14'd13064: ff_rdata <= 8'h60;
			14'd13065: ff_rdata <= 8'h00;
			14'd13066: ff_rdata <= 8'h00;
			14'd13067: ff_rdata <= 8'h00;
			14'd13068: ff_rdata <= 8'h50;
			14'd13069: ff_rdata <= 8'h69;
			14'd13070: ff_rdata <= 8'h70;
			14'd13071: ff_rdata <= 8'h65;
			14'd13072: ff_rdata <= 8'h4F;
			14'd13073: ff_rdata <= 8'h72;
			14'd13074: ff_rdata <= 8'h67;
			14'd13075: ff_rdata <= 8'h32;
			14'd13076: ff_rdata <= 8'h00;
			14'd13077: ff_rdata <= 8'h00;
			14'd13078: ff_rdata <= 8'h0C;
			14'd13079: ff_rdata <= 8'h00;
			14'd13080: ff_rdata <= 8'h00;
			14'd13081: ff_rdata <= 8'h00;
			14'd13082: ff_rdata <= 8'h00;
			14'd13083: ff_rdata <= 8'h00;
			14'd13084: ff_rdata <= 8'h34;
			14'd13085: ff_rdata <= 8'h26;
			14'd13086: ff_rdata <= 8'h50;
			14'd13087: ff_rdata <= 8'h76;
			14'd13088: ff_rdata <= 8'h30;
			14'd13089: ff_rdata <= 8'h00;
			14'd13090: ff_rdata <= 8'h00;
			14'd13091: ff_rdata <= 8'h00;
			14'd13092: ff_rdata <= 8'h30;
			14'd13093: ff_rdata <= 8'h00;
			14'd13094: ff_rdata <= 8'h30;
			14'd13095: ff_rdata <= 8'h06;
			14'd13096: ff_rdata <= 8'h80;
			14'd13097: ff_rdata <= 8'h00;
			14'd13098: ff_rdata <= 8'h00;
			14'd13099: ff_rdata <= 8'h00;
			14'd13100: ff_rdata <= 8'h50;
			14'd13101: ff_rdata <= 8'h6F;
			14'd13102: ff_rdata <= 8'h68;
			14'd13103: ff_rdata <= 8'h64;
			14'd13104: ff_rdata <= 8'h73;
			14'd13105: ff_rdata <= 8'h50;
			14'd13106: ff_rdata <= 8'h4C;
			14'd13107: ff_rdata <= 8'h41;
			14'd13108: ff_rdata <= 8'h00;
			14'd13109: ff_rdata <= 8'hED;
			14'd13110: ff_rdata <= 8'h0C;
			14'd13111: ff_rdata <= 8'h00;
			14'd13112: ff_rdata <= 8'h00;
			14'd13113: ff_rdata <= 8'h00;
			14'd13114: ff_rdata <= 8'h00;
			14'd13115: ff_rdata <= 8'h00;
			14'd13116: ff_rdata <= 8'h73;
			14'd13117: ff_rdata <= 8'h5A;
			14'd13118: ff_rdata <= 8'h99;
			14'd13119: ff_rdata <= 8'h14;
			14'd13120: ff_rdata <= 8'h60;
			14'd13121: ff_rdata <= 8'h00;
			14'd13122: ff_rdata <= 8'h00;
			14'd13123: ff_rdata <= 8'h00;
			14'd13124: ff_rdata <= 8'h33;
			14'd13125: ff_rdata <= 8'h00;
			14'd13126: ff_rdata <= 8'hF5;
			14'd13127: ff_rdata <= 8'h15;
			14'd13128: ff_rdata <= 8'h80;
			14'd13129: ff_rdata <= 8'h00;
			14'd13130: ff_rdata <= 8'h00;
			14'd13131: ff_rdata <= 8'h00;
			14'd13132: ff_rdata <= 8'h52;
			14'd13133: ff_rdata <= 8'h6F;
			14'd13134: ff_rdata <= 8'h68;
			14'd13135: ff_rdata <= 8'h64;
			14'd13136: ff_rdata <= 8'h73;
			14'd13137: ff_rdata <= 8'h50;
			14'd13138: ff_rdata <= 8'h52;
			14'd13139: ff_rdata <= 8'h41;
			14'd13140: ff_rdata <= 8'h00;
			14'd13141: ff_rdata <= 8'hED;
			14'd13142: ff_rdata <= 8'h0A;
			14'd13143: ff_rdata <= 8'h00;
			14'd13144: ff_rdata <= 8'h00;
			14'd13145: ff_rdata <= 8'h00;
			14'd13146: ff_rdata <= 8'h00;
			14'd13147: ff_rdata <= 8'h00;
			14'd13148: ff_rdata <= 8'h73;
			14'd13149: ff_rdata <= 8'h16;
			14'd13150: ff_rdata <= 8'hF9;
			14'd13151: ff_rdata <= 8'h33;
			14'd13152: ff_rdata <= 8'h60;
			14'd13153: ff_rdata <= 8'h00;
			14'd13154: ff_rdata <= 8'h00;
			14'd13155: ff_rdata <= 8'h00;
			14'd13156: ff_rdata <= 8'h13;
			14'd13157: ff_rdata <= 8'h00;
			14'd13158: ff_rdata <= 8'hF5;
			14'd13159: ff_rdata <= 8'h03;
			14'd13160: ff_rdata <= 8'h50;
			14'd13161: ff_rdata <= 8'h00;
			14'd13162: ff_rdata <= 8'h00;
			14'd13163: ff_rdata <= 8'h00;
			14'd13164: ff_rdata <= 8'h4F;
			14'd13165: ff_rdata <= 8'h72;
			14'd13166: ff_rdata <= 8'h63;
			14'd13167: ff_rdata <= 8'h68;
			14'd13168: ff_rdata <= 8'h20;
			14'd13169: ff_rdata <= 8'h4C;
			14'd13170: ff_rdata <= 8'h20;
			14'd13171: ff_rdata <= 8'h20;
			14'd13172: ff_rdata <= 8'h00;
			14'd13173: ff_rdata <= 8'h0C;
			14'd13174: ff_rdata <= 8'h0E;
			14'd13175: ff_rdata <= 8'h00;
			14'd13176: ff_rdata <= 8'h00;
			14'd13177: ff_rdata <= 8'h00;
			14'd13178: ff_rdata <= 8'h00;
			14'd13179: ff_rdata <= 8'h00;
			14'd13180: ff_rdata <= 8'h61;
			14'd13181: ff_rdata <= 8'h15;
			14'd13182: ff_rdata <= 8'h76;
			14'd13183: ff_rdata <= 8'h23;
			14'd13184: ff_rdata <= 8'h40;
			14'd13185: ff_rdata <= 8'h00;
			14'd13186: ff_rdata <= 8'h00;
			14'd13187: ff_rdata <= 8'h00;
			14'd13188: ff_rdata <= 8'h21;
			14'd13189: ff_rdata <= 8'h00;
			14'd13190: ff_rdata <= 8'h54;
			14'd13191: ff_rdata <= 8'h06;
			14'd13192: ff_rdata <= 8'h70;
			14'd13193: ff_rdata <= 8'h00;
			14'd13194: ff_rdata <= 8'h00;
			14'd13195: ff_rdata <= 8'h00;
			14'd13196: ff_rdata <= 8'h4F;
			14'd13197: ff_rdata <= 8'h72;
			14'd13198: ff_rdata <= 8'h63;
			14'd13199: ff_rdata <= 8'h68;
			14'd13200: ff_rdata <= 8'h20;
			14'd13201: ff_rdata <= 8'h52;
			14'd13202: ff_rdata <= 8'h20;
			14'd13203: ff_rdata <= 8'h20;
			14'd13204: ff_rdata <= 8'h00;
			14'd13205: ff_rdata <= 8'h00;
			14'd13206: ff_rdata <= 8'h0E;
			14'd13207: ff_rdata <= 8'h00;
			14'd13208: ff_rdata <= 8'h00;
			14'd13209: ff_rdata <= 8'h00;
			14'd13210: ff_rdata <= 8'h00;
			14'd13211: ff_rdata <= 8'h00;
			14'd13212: ff_rdata <= 8'h63;
			14'd13213: ff_rdata <= 8'h1B;
			14'd13214: ff_rdata <= 8'h75;
			14'd13215: ff_rdata <= 8'h45;
			14'd13216: ff_rdata <= 8'h60;
			14'd13217: ff_rdata <= 8'h00;
			14'd13218: ff_rdata <= 8'h00;
			14'd13219: ff_rdata <= 8'h00;
			14'd13220: ff_rdata <= 8'h70;
			14'd13221: ff_rdata <= 8'h00;
			14'd13222: ff_rdata <= 8'h4B;
			14'd13223: ff_rdata <= 8'h15;
			14'd13224: ff_rdata <= 8'h70;
			14'd13225: ff_rdata <= 8'h00;
			14'd13226: ff_rdata <= 8'h00;
			14'd13227: ff_rdata <= 8'h00;
			14'd13228: ff_rdata <= 8'h53;
			14'd13229: ff_rdata <= 8'h79;
			14'd13230: ff_rdata <= 8'h6E;
			14'd13231: ff_rdata <= 8'h56;
			14'd13232: ff_rdata <= 8'h69;
			14'd13233: ff_rdata <= 8'h6F;
			14'd13234: ff_rdata <= 8'h6C;
			14'd13235: ff_rdata <= 8'h20;
			14'd13236: ff_rdata <= 8'h00;
			14'd13237: ff_rdata <= 8'h0C;
			14'd13238: ff_rdata <= 8'h0A;
			14'd13239: ff_rdata <= 8'h00;
			14'd13240: ff_rdata <= 8'h00;
			14'd13241: ff_rdata <= 8'h00;
			14'd13242: ff_rdata <= 8'h00;
			14'd13243: ff_rdata <= 8'h00;
			14'd13244: ff_rdata <= 8'h61;
			14'd13245: ff_rdata <= 8'h0A;
			14'd13246: ff_rdata <= 8'h76;
			14'd13247: ff_rdata <= 8'h12;
			14'd13248: ff_rdata <= 8'h40;
			14'd13249: ff_rdata <= 8'h00;
			14'd13250: ff_rdata <= 8'h00;
			14'd13251: ff_rdata <= 8'h00;
			14'd13252: ff_rdata <= 8'hA1;
			14'd13253: ff_rdata <= 8'h02;
			14'd13254: ff_rdata <= 8'h54;
			14'd13255: ff_rdata <= 8'h07;
			14'd13256: ff_rdata <= 8'h80;
			14'd13257: ff_rdata <= 8'h00;
			14'd13258: ff_rdata <= 8'h00;
			14'd13259: ff_rdata <= 8'h00;
			14'd13260: ff_rdata <= 8'h53;
			14'd13261: ff_rdata <= 8'h79;
			14'd13262: ff_rdata <= 8'h6E;
			14'd13263: ff_rdata <= 8'h4F;
			14'd13264: ff_rdata <= 8'h72;
			14'd13265: ff_rdata <= 8'h67;
			14'd13266: ff_rdata <= 8'h61;
			14'd13267: ff_rdata <= 8'h6E;
			14'd13268: ff_rdata <= 8'h00;
			14'd13269: ff_rdata <= 8'hF4;
			14'd13270: ff_rdata <= 8'h0A;
			14'd13271: ff_rdata <= 8'h00;
			14'd13272: ff_rdata <= 8'h00;
			14'd13273: ff_rdata <= 8'h00;
			14'd13274: ff_rdata <= 8'h00;
			14'd13275: ff_rdata <= 8'h00;
			14'd13276: ff_rdata <= 8'h61;
			14'd13277: ff_rdata <= 8'h0D;
			14'd13278: ff_rdata <= 8'h85;
			14'd13279: ff_rdata <= 8'h14;
			14'd13280: ff_rdata <= 8'h40;
			14'd13281: ff_rdata <= 8'h00;
			14'd13282: ff_rdata <= 8'h00;
			14'd13283: ff_rdata <= 8'h00;
			14'd13284: ff_rdata <= 8'h78;
			14'd13285: ff_rdata <= 8'h08;
			14'd13286: ff_rdata <= 8'hF2;
			14'd13287: ff_rdata <= 8'h03;
			14'd13288: ff_rdata <= 8'h60;
			14'd13289: ff_rdata <= 8'h00;
			14'd13290: ff_rdata <= 8'h00;
			14'd13291: ff_rdata <= 8'h00;
			14'd13292: ff_rdata <= 8'h53;
			14'd13293: ff_rdata <= 8'h79;
			14'd13294: ff_rdata <= 8'h6E;
			14'd13295: ff_rdata <= 8'h42;
			14'd13296: ff_rdata <= 8'h72;
			14'd13297: ff_rdata <= 8'h61;
			14'd13298: ff_rdata <= 8'h73;
			14'd13299: ff_rdata <= 8'h73;
			14'd13300: ff_rdata <= 8'h00;
			14'd13301: ff_rdata <= 8'hF4;
			14'd13302: ff_rdata <= 8'h0E;
			14'd13303: ff_rdata <= 8'h00;
			14'd13304: ff_rdata <= 8'h00;
			14'd13305: ff_rdata <= 8'h00;
			14'd13306: ff_rdata <= 8'h00;
			14'd13307: ff_rdata <= 8'h00;
			14'd13308: ff_rdata <= 8'h31;
			14'd13309: ff_rdata <= 8'h15;
			14'd13310: ff_rdata <= 8'hB6;
			14'd13311: ff_rdata <= 8'h03;
			14'd13312: ff_rdata <= 8'h40;
			14'd13313: ff_rdata <= 8'h00;
			14'd13314: ff_rdata <= 8'h00;
			14'd13315: ff_rdata <= 8'h00;
			14'd13316: ff_rdata <= 8'h71;
			14'd13317: ff_rdata <= 8'h00;
			14'd13318: ff_rdata <= 8'hF9;
			14'd13319: ff_rdata <= 8'h26;
			14'd13320: ff_rdata <= 8'h60;
			14'd13321: ff_rdata <= 8'h00;
			14'd13322: ff_rdata <= 8'h00;
			14'd13323: ff_rdata <= 8'h00;
			14'd13324: ff_rdata <= 8'h54;
			14'd13325: ff_rdata <= 8'h75;
			14'd13326: ff_rdata <= 8'h62;
			14'd13327: ff_rdata <= 8'h65;
			14'd13328: ff_rdata <= 8'h20;
			14'd13329: ff_rdata <= 8'h20;
			14'd13330: ff_rdata <= 8'h20;
			14'd13331: ff_rdata <= 8'h20;
			14'd13332: ff_rdata <= 8'h00;
			14'd13333: ff_rdata <= 8'hF4;
			14'd13334: ff_rdata <= 8'h0A;
			14'd13335: ff_rdata <= 8'h00;
			14'd13336: ff_rdata <= 8'h00;
			14'd13337: ff_rdata <= 8'h00;
			14'd13338: ff_rdata <= 8'h00;
			14'd13339: ff_rdata <= 8'h00;
			14'd13340: ff_rdata <= 8'h61;
			14'd13341: ff_rdata <= 8'h0D;
			14'd13342: ff_rdata <= 8'h75;
			14'd13343: ff_rdata <= 8'h18;
			14'd13344: ff_rdata <= 8'h40;
			14'd13345: ff_rdata <= 8'h00;
			14'd13346: ff_rdata <= 8'h00;
			14'd13347: ff_rdata <= 8'h00;
			14'd13348: ff_rdata <= 8'h71;
			14'd13349: ff_rdata <= 8'h00;
			14'd13350: ff_rdata <= 8'hF2;
			14'd13351: ff_rdata <= 8'h03;
			14'd13352: ff_rdata <= 8'h60;
			14'd13353: ff_rdata <= 8'h00;
			14'd13354: ff_rdata <= 8'h00;
			14'd13355: ff_rdata <= 8'h00;
			14'd13356: ff_rdata <= 8'h53;
			14'd13357: ff_rdata <= 8'h68;
			14'd13358: ff_rdata <= 8'h61;
			14'd13359: ff_rdata <= 8'h6D;
			14'd13360: ff_rdata <= 8'h69;
			14'd13361: ff_rdata <= 8'h73;
			14'd13362: ff_rdata <= 8'h65;
			14'd13363: ff_rdata <= 8'h6E;
			14'd13364: ff_rdata <= 8'h00;
			14'd13365: ff_rdata <= 8'hED;
			14'd13366: ff_rdata <= 8'h0C;
			14'd13367: ff_rdata <= 8'h00;
			14'd13368: ff_rdata <= 8'h00;
			14'd13369: ff_rdata <= 8'h00;
			14'd13370: ff_rdata <= 8'h00;
			14'd13371: ff_rdata <= 8'h00;
			14'd13372: ff_rdata <= 8'h03;
			14'd13373: ff_rdata <= 8'h14;
			14'd13374: ff_rdata <= 8'hA7;
			14'd13375: ff_rdata <= 8'h13;
			14'd13376: ff_rdata <= 8'h50;
			14'd13377: ff_rdata <= 8'h00;
			14'd13378: ff_rdata <= 8'h00;
			14'd13379: ff_rdata <= 8'h00;
			14'd13380: ff_rdata <= 8'h0C;
			14'd13381: ff_rdata <= 8'h03;
			14'd13382: ff_rdata <= 8'hFC;
			14'd13383: ff_rdata <= 8'h15;
			14'd13384: ff_rdata <= 8'h60;
			14'd13385: ff_rdata <= 8'h00;
			14'd13386: ff_rdata <= 8'h00;
			14'd13387: ff_rdata <= 8'h00;
			14'd13388: ff_rdata <= 8'h4D;
			14'd13389: ff_rdata <= 8'h61;
			14'd13390: ff_rdata <= 8'h67;
			14'd13391: ff_rdata <= 8'h69;
			14'd13392: ff_rdata <= 8'h63;
			14'd13393: ff_rdata <= 8'h61;
			14'd13394: ff_rdata <= 8'h6C;
			14'd13395: ff_rdata <= 8'h20;
			14'd13396: ff_rdata <= 8'h00;
			14'd13397: ff_rdata <= 8'hF4;
			14'd13398: ff_rdata <= 8'h06;
			14'd13399: ff_rdata <= 8'h00;
			14'd13400: ff_rdata <= 8'h00;
			14'd13401: ff_rdata <= 8'h00;
			14'd13402: ff_rdata <= 8'h00;
			14'd13403: ff_rdata <= 8'h00;
			14'd13404: ff_rdata <= 8'h13;
			14'd13405: ff_rdata <= 8'h80;
			14'd13406: ff_rdata <= 8'h20;
			14'd13407: ff_rdata <= 8'h03;
			14'd13408: ff_rdata <= 8'h60;
			14'd13409: ff_rdata <= 8'h00;
			14'd13410: ff_rdata <= 8'h00;
			14'd13411: ff_rdata <= 8'h00;
			14'd13412: ff_rdata <= 8'h32;
			14'd13413: ff_rdata <= 8'h00;
			14'd13414: ff_rdata <= 8'h85;
			14'd13415: ff_rdata <= 8'hAF;
			14'd13416: ff_rdata <= 8'h40;
			14'd13417: ff_rdata <= 8'h00;
			14'd13418: ff_rdata <= 8'h00;
			14'd13419: ff_rdata <= 8'h00;
			14'd13420: ff_rdata <= 8'h48;
			14'd13421: ff_rdata <= 8'h75;
			14'd13422: ff_rdata <= 8'h77;
			14'd13423: ff_rdata <= 8'h61;
			14'd13424: ff_rdata <= 8'h77;
			14'd13425: ff_rdata <= 8'h61;
			14'd13426: ff_rdata <= 8'h20;
			14'd13427: ff_rdata <= 8'h20;
			14'd13428: ff_rdata <= 8'h00;
			14'd13429: ff_rdata <= 8'h00;
			14'd13430: ff_rdata <= 8'h0A;
			14'd13431: ff_rdata <= 8'h00;
			14'd13432: ff_rdata <= 8'h00;
			14'd13433: ff_rdata <= 8'h00;
			14'd13434: ff_rdata <= 8'h00;
			14'd13435: ff_rdata <= 8'h00;
			14'd13436: ff_rdata <= 8'hF1;
			14'd13437: ff_rdata <= 8'h17;
			14'd13438: ff_rdata <= 8'h23;
			14'd13439: ff_rdata <= 8'h14;
			14'd13440: ff_rdata <= 8'h20;
			14'd13441: ff_rdata <= 8'h00;
			14'd13442: ff_rdata <= 8'h00;
			14'd13443: ff_rdata <= 8'h00;
			14'd13444: ff_rdata <= 8'h31;
			14'd13445: ff_rdata <= 8'h00;
			14'd13446: ff_rdata <= 8'h40;
			14'd13447: ff_rdata <= 8'h09;
			14'd13448: ff_rdata <= 8'h80;
			14'd13449: ff_rdata <= 8'h00;
			14'd13450: ff_rdata <= 8'h00;
			14'd13451: ff_rdata <= 8'h00;
			14'd13452: ff_rdata <= 8'h57;
			14'd13453: ff_rdata <= 8'h6E;
			14'd13454: ff_rdata <= 8'h64;
			14'd13455: ff_rdata <= 8'h65;
			14'd13456: ff_rdata <= 8'h72;
			14'd13457: ff_rdata <= 8'h46;
			14'd13458: ff_rdata <= 8'h6C;
			14'd13459: ff_rdata <= 8'h74;
			14'd13460: ff_rdata <= 8'h00;
			14'd13461: ff_rdata <= 8'h00;
			14'd13462: ff_rdata <= 8'hEE;
			14'd13463: ff_rdata <= 8'h00;
			14'd13464: ff_rdata <= 8'h00;
			14'd13465: ff_rdata <= 8'h00;
			14'd13466: ff_rdata <= 8'h00;
			14'd13467: ff_rdata <= 8'h00;
			14'd13468: ff_rdata <= 8'hF0;
			14'd13469: ff_rdata <= 8'h17;
			14'd13470: ff_rdata <= 8'h5A;
			14'd13471: ff_rdata <= 8'h06;
			14'd13472: ff_rdata <= 8'h40;
			14'd13473: ff_rdata <= 8'h00;
			14'd13474: ff_rdata <= 8'h00;
			14'd13475: ff_rdata <= 8'h00;
			14'd13476: ff_rdata <= 8'h74;
			14'd13477: ff_rdata <= 8'h40;
			14'd13478: ff_rdata <= 8'h43;
			14'd13479: ff_rdata <= 8'hFC;
			14'd13480: ff_rdata <= 8'h80;
			14'd13481: ff_rdata <= 8'h00;
			14'd13482: ff_rdata <= 8'h00;
			14'd13483: ff_rdata <= 8'h00;
			14'd13484: ff_rdata <= 8'h48;
			14'd13485: ff_rdata <= 8'h61;
			14'd13486: ff_rdata <= 8'h72;
			14'd13487: ff_rdata <= 8'h64;
			14'd13488: ff_rdata <= 8'h72;
			14'd13489: ff_rdata <= 8'h6F;
			14'd13490: ff_rdata <= 8'h63;
			14'd13491: ff_rdata <= 8'h6B;
			14'd13492: ff_rdata <= 8'h00;
			14'd13493: ff_rdata <= 8'h00;
			14'd13494: ff_rdata <= 8'h6C;
			14'd13495: ff_rdata <= 8'h00;
			14'd13496: ff_rdata <= 8'h00;
			14'd13497: ff_rdata <= 8'h00;
			14'd13498: ff_rdata <= 8'h00;
			14'd13499: ff_rdata <= 8'h00;
			14'd13500: ff_rdata <= 8'h20;
			14'd13501: ff_rdata <= 8'h0D;
			14'd13502: ff_rdata <= 8'hC1;
			14'd13503: ff_rdata <= 8'h56;
			14'd13504: ff_rdata <= 8'h20;
			14'd13505: ff_rdata <= 8'h00;
			14'd13506: ff_rdata <= 8'h00;
			14'd13507: ff_rdata <= 8'h00;
			14'd13508: ff_rdata <= 8'h71;
			14'd13509: ff_rdata <= 8'h02;
			14'd13510: ff_rdata <= 8'hD5;
			14'd13511: ff_rdata <= 8'h06;
			14'd13512: ff_rdata <= 8'h60;
			14'd13513: ff_rdata <= 8'h00;
			14'd13514: ff_rdata <= 8'h00;
			14'd13515: ff_rdata <= 8'h00;
			14'd13516: ff_rdata <= 8'h4D;
			14'd13517: ff_rdata <= 8'h61;
			14'd13518: ff_rdata <= 8'h63;
			14'd13519: ff_rdata <= 8'h68;
			14'd13520: ff_rdata <= 8'h69;
			14'd13521: ff_rdata <= 8'h6E;
			14'd13522: ff_rdata <= 8'h65;
			14'd13523: ff_rdata <= 8'h20;
			14'd13524: ff_rdata <= 8'h00;
			14'd13525: ff_rdata <= 8'hF4;
			14'd13526: ff_rdata <= 8'h0C;
			14'd13527: ff_rdata <= 8'h00;
			14'd13528: ff_rdata <= 8'h00;
			14'd13529: ff_rdata <= 8'h00;
			14'd13530: ff_rdata <= 8'h00;
			14'd13531: ff_rdata <= 8'h00;
			14'd13532: ff_rdata <= 8'h30;
			14'd13533: ff_rdata <= 8'h06;
			14'd13534: ff_rdata <= 8'h40;
			14'd13535: ff_rdata <= 8'h04;
			14'd13536: ff_rdata <= 8'h80;
			14'd13537: ff_rdata <= 8'h00;
			14'd13538: ff_rdata <= 8'h00;
			14'd13539: ff_rdata <= 8'h00;
			14'd13540: ff_rdata <= 8'h32;
			14'd13541: ff_rdata <= 8'h00;
			14'd13542: ff_rdata <= 8'h40;
			14'd13543: ff_rdata <= 8'h74;
			14'd13544: ff_rdata <= 8'h30;
			14'd13545: ff_rdata <= 8'h00;
			14'd13546: ff_rdata <= 8'h00;
			14'd13547: ff_rdata <= 8'h00;
			14'd13548: ff_rdata <= 8'h4D;
			14'd13549: ff_rdata <= 8'h61;
			14'd13550: ff_rdata <= 8'h63;
			14'd13551: ff_rdata <= 8'h68;
			14'd13552: ff_rdata <= 8'h69;
			14'd13553: ff_rdata <= 8'h6E;
			14'd13554: ff_rdata <= 8'h65;
			14'd13555: ff_rdata <= 8'h56;
			14'd13556: ff_rdata <= 8'h00;
			14'd13557: ff_rdata <= 8'hF4;
			14'd13558: ff_rdata <= 8'h06;
			14'd13559: ff_rdata <= 8'h00;
			14'd13560: ff_rdata <= 8'h00;
			14'd13561: ff_rdata <= 8'h00;
			14'd13562: ff_rdata <= 8'h00;
			14'd13563: ff_rdata <= 8'h00;
			14'd13564: ff_rdata <= 8'h30;
			14'd13565: ff_rdata <= 8'h03;
			14'd13566: ff_rdata <= 8'h40;
			14'd13567: ff_rdata <= 8'h04;
			14'd13568: ff_rdata <= 8'h80;
			14'd13569: ff_rdata <= 8'h00;
			14'd13570: ff_rdata <= 8'h00;
			14'd13571: ff_rdata <= 8'h00;
			14'd13572: ff_rdata <= 8'h32;
			14'd13573: ff_rdata <= 8'h00;
			14'd13574: ff_rdata <= 8'h40;
			14'd13575: ff_rdata <= 8'h74;
			14'd13576: ff_rdata <= 8'h30;
			14'd13577: ff_rdata <= 8'h00;
			14'd13578: ff_rdata <= 8'h00;
			14'd13579: ff_rdata <= 8'h00;
			14'd13580: ff_rdata <= 8'h43;
			14'd13581: ff_rdata <= 8'h6F;
			14'd13582: ff_rdata <= 8'h6D;
			14'd13583: ff_rdata <= 8'h69;
			14'd13584: ff_rdata <= 8'h63;
			14'd13585: ff_rdata <= 8'h20;
			14'd13586: ff_rdata <= 8'h20;
			14'd13587: ff_rdata <= 8'h20;
			14'd13588: ff_rdata <= 8'h00;
			14'd13589: ff_rdata <= 8'hF4;
			14'd13590: ff_rdata <= 8'h0E;
			14'd13591: ff_rdata <= 8'h00;
			14'd13592: ff_rdata <= 8'h00;
			14'd13593: ff_rdata <= 8'h00;
			14'd13594: ff_rdata <= 8'h00;
			14'd13595: ff_rdata <= 8'h00;
			14'd13596: ff_rdata <= 8'h01;
			14'd13597: ff_rdata <= 8'h0D;
			14'd13598: ff_rdata <= 8'h78;
			14'd13599: ff_rdata <= 8'h7F;
			14'd13600: ff_rdata <= 8'h40;
			14'd13601: ff_rdata <= 8'h00;
			14'd13602: ff_rdata <= 8'h00;
			14'd13603: ff_rdata <= 8'h00;
			14'd13604: ff_rdata <= 8'h08;
			14'd13605: ff_rdata <= 8'h00;
			14'd13606: ff_rdata <= 8'hF8;
			14'd13607: ff_rdata <= 8'hF9;
			14'd13608: ff_rdata <= 8'h00;
			14'd13609: ff_rdata <= 8'h00;
			14'd13610: ff_rdata <= 8'h00;
			14'd13611: ff_rdata <= 8'h00;
			14'd13612: ff_rdata <= 8'h53;
			14'd13613: ff_rdata <= 8'h45;
			14'd13614: ff_rdata <= 8'h5F;
			14'd13615: ff_rdata <= 8'h43;
			14'd13616: ff_rdata <= 8'h6F;
			14'd13617: ff_rdata <= 8'h6D;
			14'd13618: ff_rdata <= 8'h69;
			14'd13619: ff_rdata <= 8'h63;
			14'd13620: ff_rdata <= 8'h00;
			14'd13621: ff_rdata <= 8'hE8;
			14'd13622: ff_rdata <= 8'h6A;
			14'd13623: ff_rdata <= 8'h00;
			14'd13624: ff_rdata <= 8'h00;
			14'd13625: ff_rdata <= 8'h00;
			14'd13626: ff_rdata <= 8'h00;
			14'd13627: ff_rdata <= 8'h00;
			14'd13628: ff_rdata <= 8'hC8;
			14'd13629: ff_rdata <= 8'h0B;
			14'd13630: ff_rdata <= 8'h76;
			14'd13631: ff_rdata <= 8'h11;
			14'd13632: ff_rdata <= 8'h40;
			14'd13633: ff_rdata <= 8'h00;
			14'd13634: ff_rdata <= 8'h00;
			14'd13635: ff_rdata <= 8'h00;
			14'd13636: ff_rdata <= 8'hC0;
			14'd13637: ff_rdata <= 8'h00;
			14'd13638: ff_rdata <= 8'hF7;
			14'd13639: ff_rdata <= 8'hF9;
			14'd13640: ff_rdata <= 8'h00;
			14'd13641: ff_rdata <= 8'h00;
			14'd13642: ff_rdata <= 8'h00;
			14'd13643: ff_rdata <= 8'h00;
			14'd13644: ff_rdata <= 8'h53;
			14'd13645: ff_rdata <= 8'h45;
			14'd13646: ff_rdata <= 8'h5F;
			14'd13647: ff_rdata <= 8'h4C;
			14'd13648: ff_rdata <= 8'h61;
			14'd13649: ff_rdata <= 8'h73;
			14'd13650: ff_rdata <= 8'h65;
			14'd13651: ff_rdata <= 8'h72;
			14'd13652: ff_rdata <= 8'h00;
			14'd13653: ff_rdata <= 8'h30;
			14'd13654: ff_rdata <= 8'h6E;
			14'd13655: ff_rdata <= 8'h00;
			14'd13656: ff_rdata <= 8'h00;
			14'd13657: ff_rdata <= 8'h00;
			14'd13658: ff_rdata <= 8'h00;
			14'd13659: ff_rdata <= 8'h00;
			14'd13660: ff_rdata <= 8'h49;
			14'd13661: ff_rdata <= 8'h0B;
			14'd13662: ff_rdata <= 8'hB4;
			14'd13663: ff_rdata <= 8'hFF;
			14'd13664: ff_rdata <= 8'h20;
			14'd13665: ff_rdata <= 8'h00;
			14'd13666: ff_rdata <= 8'h00;
			14'd13667: ff_rdata <= 8'h00;
			14'd13668: ff_rdata <= 8'h40;
			14'd13669: ff_rdata <= 8'h00;
			14'd13670: ff_rdata <= 8'hF9;
			14'd13671: ff_rdata <= 8'h05;
			14'd13672: ff_rdata <= 8'h60;
			14'd13673: ff_rdata <= 8'h00;
			14'd13674: ff_rdata <= 8'h00;
			14'd13675: ff_rdata <= 8'h00;
			14'd13676: ff_rdata <= 8'h53;
			14'd13677: ff_rdata <= 8'h45;
			14'd13678: ff_rdata <= 8'h5F;
			14'd13679: ff_rdata <= 8'h4E;
			14'd13680: ff_rdata <= 8'h6F;
			14'd13681: ff_rdata <= 8'h69;
			14'd13682: ff_rdata <= 8'h73;
			14'd13683: ff_rdata <= 8'h65;
			14'd13684: ff_rdata <= 8'h00;
			14'd13685: ff_rdata <= 8'h24;
			14'd13686: ff_rdata <= 8'hAC;
			14'd13687: ff_rdata <= 8'h00;
			14'd13688: ff_rdata <= 8'h00;
			14'd13689: ff_rdata <= 8'h00;
			14'd13690: ff_rdata <= 8'h00;
			14'd13691: ff_rdata <= 8'h00;
			14'd13692: ff_rdata <= 8'hCD;
			14'd13693: ff_rdata <= 8'h0C;
			14'd13694: ff_rdata <= 8'hA2;
			14'd13695: ff_rdata <= 8'h00;
			14'd13696: ff_rdata <= 8'h80;
			14'd13697: ff_rdata <= 8'h00;
			14'd13698: ff_rdata <= 8'h00;
			14'd13699: ff_rdata <= 8'h00;
			14'd13700: ff_rdata <= 8'h42;
			14'd13701: ff_rdata <= 8'h00;
			14'd13702: ff_rdata <= 8'hF0;
			14'd13703: ff_rdata <= 8'h01;
			14'd13704: ff_rdata <= 8'h80;
			14'd13705: ff_rdata <= 8'h00;
			14'd13706: ff_rdata <= 8'h00;
			14'd13707: ff_rdata <= 8'h00;
			14'd13708: ff_rdata <= 8'h53;
			14'd13709: ff_rdata <= 8'h45;
			14'd13710: ff_rdata <= 8'h5F;
			14'd13711: ff_rdata <= 8'h53;
			14'd13712: ff_rdata <= 8'h74;
			14'd13713: ff_rdata <= 8'h61;
			14'd13714: ff_rdata <= 8'h72;
			14'd13715: ff_rdata <= 8'h20;
			14'd13716: ff_rdata <= 8'h00;
			14'd13717: ff_rdata <= 8'h00;
			14'd13718: ff_rdata <= 8'h6E;
			14'd13719: ff_rdata <= 8'h00;
			14'd13720: ff_rdata <= 8'h00;
			14'd13721: ff_rdata <= 8'h00;
			14'd13722: ff_rdata <= 8'h00;
			14'd13723: ff_rdata <= 8'h00;
			14'd13724: ff_rdata <= 8'h51;
			14'd13725: ff_rdata <= 8'h13;
			14'd13726: ff_rdata <= 8'h13;
			14'd13727: ff_rdata <= 8'h42;
			14'd13728: ff_rdata <= 8'h40;
			14'd13729: ff_rdata <= 8'h00;
			14'd13730: ff_rdata <= 8'h00;
			14'd13731: ff_rdata <= 8'h00;
			14'd13732: ff_rdata <= 8'h42;
			14'd13733: ff_rdata <= 8'h00;
			14'd13734: ff_rdata <= 8'h10;
			14'd13735: ff_rdata <= 8'h01;
			14'd13736: ff_rdata <= 8'h50;
			14'd13737: ff_rdata <= 8'h00;
			14'd13738: ff_rdata <= 8'h00;
			14'd13739: ff_rdata <= 8'h00;
			14'd13740: ff_rdata <= 8'h53;
			14'd13741: ff_rdata <= 8'h45;
			14'd13742: ff_rdata <= 8'h5F;
			14'd13743: ff_rdata <= 8'h53;
			14'd13744: ff_rdata <= 8'h74;
			14'd13745: ff_rdata <= 8'h61;
			14'd13746: ff_rdata <= 8'h72;
			14'd13747: ff_rdata <= 8'h32;
			14'd13748: ff_rdata <= 8'h00;
			14'd13749: ff_rdata <= 8'h24;
			14'd13750: ff_rdata <= 8'h6E;
			14'd13751: ff_rdata <= 8'h00;
			14'd13752: ff_rdata <= 8'h00;
			14'd13753: ff_rdata <= 8'h00;
			14'd13754: ff_rdata <= 8'h00;
			14'd13755: ff_rdata <= 8'h00;
			14'd13756: ff_rdata <= 8'h51;
			14'd13757: ff_rdata <= 8'h13;
			14'd13758: ff_rdata <= 8'h13;
			14'd13759: ff_rdata <= 8'h42;
			14'd13760: ff_rdata <= 8'h40;
			14'd13761: ff_rdata <= 8'h00;
			14'd13762: ff_rdata <= 8'h00;
			14'd13763: ff_rdata <= 8'h00;
			14'd13764: ff_rdata <= 8'h42;
			14'd13765: ff_rdata <= 8'h00;
			14'd13766: ff_rdata <= 8'h10;
			14'd13767: ff_rdata <= 8'h01;
			14'd13768: ff_rdata <= 8'h50;
			14'd13769: ff_rdata <= 8'h00;
			14'd13770: ff_rdata <= 8'h00;
			14'd13771: ff_rdata <= 8'h00;
			14'd13772: ff_rdata <= 8'h45;
			14'd13773: ff_rdata <= 8'h6E;
			14'd13774: ff_rdata <= 8'h67;
			14'd13775: ff_rdata <= 8'h69;
			14'd13776: ff_rdata <= 8'h6E;
			14'd13777: ff_rdata <= 8'h65;
			14'd13778: ff_rdata <= 8'h20;
			14'd13779: ff_rdata <= 8'h32;
			14'd13780: ff_rdata <= 8'h00;
			14'd13781: ff_rdata <= 8'hE8;
			14'd13782: ff_rdata <= 8'h0C;
			14'd13783: ff_rdata <= 8'h00;
			14'd13784: ff_rdata <= 8'h00;
			14'd13785: ff_rdata <= 8'h00;
			14'd13786: ff_rdata <= 8'h00;
			14'd13787: ff_rdata <= 8'h00;
			14'd13788: ff_rdata <= 8'h30;
			14'd13789: ff_rdata <= 8'h12;
			14'd13790: ff_rdata <= 8'h23;
			14'd13791: ff_rdata <= 8'h26;
			14'd13792: ff_rdata <= 8'h40;
			14'd13793: ff_rdata <= 8'h00;
			14'd13794: ff_rdata <= 8'h00;
			14'd13795: ff_rdata <= 8'h00;
			14'd13796: ff_rdata <= 8'h34;
			14'd13797: ff_rdata <= 8'h07;
			14'd13798: ff_rdata <= 8'h70;
			14'd13799: ff_rdata <= 8'h02;
			14'd13800: ff_rdata <= 8'h50;
			14'd13801: ff_rdata <= 8'h00;
			14'd13802: ff_rdata <= 8'h00;
			14'd13803: ff_rdata <= 8'h00;
			14'd13804: ff_rdata <= 8'h53;
			14'd13805: ff_rdata <= 8'h69;
			14'd13806: ff_rdata <= 8'h6C;
			14'd13807: ff_rdata <= 8'h65;
			14'd13808: ff_rdata <= 8'h6E;
			14'd13809: ff_rdata <= 8'h63;
			14'd13810: ff_rdata <= 8'h65;
			14'd13811: ff_rdata <= 8'h20;
			14'd13812: ff_rdata <= 8'h00;
			14'd13813: ff_rdata <= 8'h00;
			14'd13814: ff_rdata <= 8'h00;
			14'd13815: ff_rdata <= 8'h00;
			14'd13816: ff_rdata <= 8'h00;
			14'd13817: ff_rdata <= 8'h00;
			14'd13818: ff_rdata <= 8'h00;
			14'd13819: ff_rdata <= 8'h00;
			14'd13820: ff_rdata <= 8'h00;
			14'd13821: ff_rdata <= 8'hFF;
			14'd13822: ff_rdata <= 8'h00;
			14'd13823: ff_rdata <= 8'hFF;
			14'd13824: ff_rdata <= 8'h00;
			14'd13825: ff_rdata <= 8'h00;
			14'd13826: ff_rdata <= 8'h00;
			14'd13827: ff_rdata <= 8'h00;
			14'd13828: ff_rdata <= 8'h00;
			14'd13829: ff_rdata <= 8'hFF;
			14'd13830: ff_rdata <= 8'h00;
			14'd13831: ff_rdata <= 8'hFF;
			14'd13832: ff_rdata <= 8'h00;
			14'd13833: ff_rdata <= 8'h00;
			14'd13834: ff_rdata <= 8'h00;
			14'd13835: ff_rdata <= 8'h00;
			14'd13836: ff_rdata <= 8'hFF;
			14'd13837: ff_rdata <= 8'hFF;
			14'd13838: ff_rdata <= 8'hFF;
			14'd13839: ff_rdata <= 8'hFF;
			14'd13840: ff_rdata <= 8'hFF;
			14'd13841: ff_rdata <= 8'hFF;
			14'd13842: ff_rdata <= 8'hFF;
			14'd13843: ff_rdata <= 8'hFF;
			14'd13844: ff_rdata <= 8'hFF;
			14'd13845: ff_rdata <= 8'hFF;
			14'd13846: ff_rdata <= 8'hFF;
			14'd13847: ff_rdata <= 8'hFF;
			14'd13848: ff_rdata <= 8'hFF;
			14'd13849: ff_rdata <= 8'hFF;
			14'd13850: ff_rdata <= 8'hFF;
			14'd13851: ff_rdata <= 8'hFF;
			14'd13852: ff_rdata <= 8'hFF;
			14'd13853: ff_rdata <= 8'hFF;
			14'd13854: ff_rdata <= 8'hFF;
			14'd13855: ff_rdata <= 8'hFF;
			14'd13856: ff_rdata <= 8'hFF;
			14'd13857: ff_rdata <= 8'hFF;
			14'd13858: ff_rdata <= 8'hFF;
			14'd13859: ff_rdata <= 8'hFF;
			14'd13860: ff_rdata <= 8'hFF;
			14'd13861: ff_rdata <= 8'hFF;
			14'd13862: ff_rdata <= 8'hFF;
			14'd13863: ff_rdata <= 8'hFF;
			14'd13864: ff_rdata <= 8'hFF;
			14'd13865: ff_rdata <= 8'hFF;
			14'd13866: ff_rdata <= 8'hFF;
			14'd13867: ff_rdata <= 8'hFF;
			14'd13868: ff_rdata <= 8'hFF;
			14'd13869: ff_rdata <= 8'hFF;
			14'd13870: ff_rdata <= 8'hFF;
			14'd13871: ff_rdata <= 8'hFF;
			14'd13872: ff_rdata <= 8'hFF;
			14'd13873: ff_rdata <= 8'hFF;
			14'd13874: ff_rdata <= 8'hFF;
			14'd13875: ff_rdata <= 8'hFF;
			14'd13876: ff_rdata <= 8'hFF;
			14'd13877: ff_rdata <= 8'hFF;
			14'd13878: ff_rdata <= 8'hFF;
			14'd13879: ff_rdata <= 8'hFF;
			14'd13880: ff_rdata <= 8'hFF;
			14'd13881: ff_rdata <= 8'hFF;
			14'd13882: ff_rdata <= 8'hFF;
			14'd13883: ff_rdata <= 8'hFF;
			14'd13884: ff_rdata <= 8'hFF;
			14'd13885: ff_rdata <= 8'hFF;
			14'd13886: ff_rdata <= 8'hFF;
			14'd13887: ff_rdata <= 8'hFF;
			14'd13888: ff_rdata <= 8'hFF;
			14'd13889: ff_rdata <= 8'hFF;
			14'd13890: ff_rdata <= 8'hFF;
			14'd13891: ff_rdata <= 8'hFF;
			14'd13892: ff_rdata <= 8'hFF;
			14'd13893: ff_rdata <= 8'hFF;
			14'd13894: ff_rdata <= 8'hFF;
			14'd13895: ff_rdata <= 8'hFF;
			14'd13896: ff_rdata <= 8'hFF;
			14'd13897: ff_rdata <= 8'hFF;
			14'd13898: ff_rdata <= 8'hFF;
			14'd13899: ff_rdata <= 8'hFF;
			14'd13900: ff_rdata <= 8'hFF;
			14'd13901: ff_rdata <= 8'hFF;
			14'd13902: ff_rdata <= 8'hFF;
			14'd13903: ff_rdata <= 8'hFF;
			14'd13904: ff_rdata <= 8'hFF;
			14'd13905: ff_rdata <= 8'hFF;
			14'd13906: ff_rdata <= 8'hFF;
			14'd13907: ff_rdata <= 8'hFF;
			14'd13908: ff_rdata <= 8'hFF;
			14'd13909: ff_rdata <= 8'hFF;
			14'd13910: ff_rdata <= 8'hFF;
			14'd13911: ff_rdata <= 8'hFF;
			14'd13912: ff_rdata <= 8'hFF;
			14'd13913: ff_rdata <= 8'hFF;
			14'd13914: ff_rdata <= 8'hFF;
			14'd13915: ff_rdata <= 8'hFF;
			14'd13916: ff_rdata <= 8'hFF;
			14'd13917: ff_rdata <= 8'hFF;
			14'd13918: ff_rdata <= 8'hFF;
			14'd13919: ff_rdata <= 8'hFF;
			14'd13920: ff_rdata <= 8'hFF;
			14'd13921: ff_rdata <= 8'hFF;
			14'd13922: ff_rdata <= 8'hFF;
			14'd13923: ff_rdata <= 8'hFF;
			14'd13924: ff_rdata <= 8'hFF;
			14'd13925: ff_rdata <= 8'hFF;
			14'd13926: ff_rdata <= 8'hFF;
			14'd13927: ff_rdata <= 8'hFF;
			14'd13928: ff_rdata <= 8'hFF;
			14'd13929: ff_rdata <= 8'hFF;
			14'd13930: ff_rdata <= 8'hFF;
			14'd13931: ff_rdata <= 8'hFF;
			14'd13932: ff_rdata <= 8'hFF;
			14'd13933: ff_rdata <= 8'hFF;
			14'd13934: ff_rdata <= 8'hFF;
			14'd13935: ff_rdata <= 8'hFF;
			14'd13936: ff_rdata <= 8'hFF;
			14'd13937: ff_rdata <= 8'hFF;
			14'd13938: ff_rdata <= 8'hFF;
			14'd13939: ff_rdata <= 8'hFF;
			14'd13940: ff_rdata <= 8'hFF;
			14'd13941: ff_rdata <= 8'hFF;
			14'd13942: ff_rdata <= 8'hFF;
			14'd13943: ff_rdata <= 8'hFF;
			14'd13944: ff_rdata <= 8'hFF;
			14'd13945: ff_rdata <= 8'hFF;
			14'd13946: ff_rdata <= 8'hFF;
			14'd13947: ff_rdata <= 8'hFF;
			14'd13948: ff_rdata <= 8'hFF;
			14'd13949: ff_rdata <= 8'hFF;
			14'd13950: ff_rdata <= 8'hFF;
			14'd13951: ff_rdata <= 8'hFF;
			14'd13952: ff_rdata <= 8'hFF;
			14'd13953: ff_rdata <= 8'hFF;
			14'd13954: ff_rdata <= 8'hFF;
			14'd13955: ff_rdata <= 8'hFF;
			14'd13956: ff_rdata <= 8'hFF;
			14'd13957: ff_rdata <= 8'hFF;
			14'd13958: ff_rdata <= 8'hFF;
			14'd13959: ff_rdata <= 8'hFF;
			14'd13960: ff_rdata <= 8'hFF;
			14'd13961: ff_rdata <= 8'hFF;
			14'd13962: ff_rdata <= 8'hFF;
			14'd13963: ff_rdata <= 8'hFF;
			14'd13964: ff_rdata <= 8'hFF;
			14'd13965: ff_rdata <= 8'hFF;
			14'd13966: ff_rdata <= 8'hFF;
			14'd13967: ff_rdata <= 8'hFF;
			14'd13968: ff_rdata <= 8'hFF;
			14'd13969: ff_rdata <= 8'hFF;
			14'd13970: ff_rdata <= 8'hFF;
			14'd13971: ff_rdata <= 8'hFF;
			14'd13972: ff_rdata <= 8'hFF;
			14'd13973: ff_rdata <= 8'hFF;
			14'd13974: ff_rdata <= 8'hFF;
			14'd13975: ff_rdata <= 8'hFF;
			14'd13976: ff_rdata <= 8'hFF;
			14'd13977: ff_rdata <= 8'hFF;
			14'd13978: ff_rdata <= 8'hFF;
			14'd13979: ff_rdata <= 8'hFF;
			14'd13980: ff_rdata <= 8'hFF;
			14'd13981: ff_rdata <= 8'hFF;
			14'd13982: ff_rdata <= 8'hFF;
			14'd13983: ff_rdata <= 8'hFF;
			14'd13984: ff_rdata <= 8'hFF;
			14'd13985: ff_rdata <= 8'hFF;
			14'd13986: ff_rdata <= 8'hFF;
			14'd13987: ff_rdata <= 8'hFF;
			14'd13988: ff_rdata <= 8'hFF;
			14'd13989: ff_rdata <= 8'hFF;
			14'd13990: ff_rdata <= 8'hFF;
			14'd13991: ff_rdata <= 8'hFF;
			14'd13992: ff_rdata <= 8'hFF;
			14'd13993: ff_rdata <= 8'hFF;
			14'd13994: ff_rdata <= 8'hFF;
			14'd13995: ff_rdata <= 8'hFF;
			14'd13996: ff_rdata <= 8'hFF;
			14'd13997: ff_rdata <= 8'hFF;
			14'd13998: ff_rdata <= 8'hFF;
			14'd13999: ff_rdata <= 8'hFF;
			14'd14000: ff_rdata <= 8'hFF;
			14'd14001: ff_rdata <= 8'hFF;
			14'd14002: ff_rdata <= 8'hFF;
			14'd14003: ff_rdata <= 8'hFF;
			14'd14004: ff_rdata <= 8'hFF;
			14'd14005: ff_rdata <= 8'hFF;
			14'd14006: ff_rdata <= 8'hFF;
			14'd14007: ff_rdata <= 8'hFF;
			14'd14008: ff_rdata <= 8'hFF;
			14'd14009: ff_rdata <= 8'hFF;
			14'd14010: ff_rdata <= 8'hFF;
			14'd14011: ff_rdata <= 8'hFF;
			14'd14012: ff_rdata <= 8'hFF;
			14'd14013: ff_rdata <= 8'hFF;
			14'd14014: ff_rdata <= 8'hFF;
			14'd14015: ff_rdata <= 8'hFF;
			14'd14016: ff_rdata <= 8'hFF;
			14'd14017: ff_rdata <= 8'hFF;
			14'd14018: ff_rdata <= 8'hFF;
			14'd14019: ff_rdata <= 8'hFF;
			14'd14020: ff_rdata <= 8'hFF;
			14'd14021: ff_rdata <= 8'hFF;
			14'd14022: ff_rdata <= 8'hFF;
			14'd14023: ff_rdata <= 8'hFF;
			14'd14024: ff_rdata <= 8'hFF;
			14'd14025: ff_rdata <= 8'hFF;
			14'd14026: ff_rdata <= 8'hFF;
			14'd14027: ff_rdata <= 8'hFF;
			14'd14028: ff_rdata <= 8'hFF;
			14'd14029: ff_rdata <= 8'hFF;
			14'd14030: ff_rdata <= 8'hFF;
			14'd14031: ff_rdata <= 8'hFF;
			14'd14032: ff_rdata <= 8'hFF;
			14'd14033: ff_rdata <= 8'hFF;
			14'd14034: ff_rdata <= 8'hFF;
			14'd14035: ff_rdata <= 8'hFF;
			14'd14036: ff_rdata <= 8'hFF;
			14'd14037: ff_rdata <= 8'hFF;
			14'd14038: ff_rdata <= 8'hFF;
			14'd14039: ff_rdata <= 8'hFF;
			14'd14040: ff_rdata <= 8'hFF;
			14'd14041: ff_rdata <= 8'hFF;
			14'd14042: ff_rdata <= 8'hFF;
			14'd14043: ff_rdata <= 8'hFF;
			14'd14044: ff_rdata <= 8'hFF;
			14'd14045: ff_rdata <= 8'hFF;
			14'd14046: ff_rdata <= 8'hFF;
			14'd14047: ff_rdata <= 8'hFF;
			14'd14048: ff_rdata <= 8'hFF;
			14'd14049: ff_rdata <= 8'hFF;
			14'd14050: ff_rdata <= 8'hFF;
			14'd14051: ff_rdata <= 8'hFF;
			14'd14052: ff_rdata <= 8'hFF;
			14'd14053: ff_rdata <= 8'hFF;
			14'd14054: ff_rdata <= 8'hFF;
			14'd14055: ff_rdata <= 8'hFF;
			14'd14056: ff_rdata <= 8'hFF;
			14'd14057: ff_rdata <= 8'hFF;
			14'd14058: ff_rdata <= 8'hFF;
			14'd14059: ff_rdata <= 8'hFF;
			14'd14060: ff_rdata <= 8'hFF;
			14'd14061: ff_rdata <= 8'hFF;
			14'd14062: ff_rdata <= 8'hFF;
			14'd14063: ff_rdata <= 8'hFF;
			14'd14064: ff_rdata <= 8'hFF;
			14'd14065: ff_rdata <= 8'hFF;
			14'd14066: ff_rdata <= 8'hFF;
			14'd14067: ff_rdata <= 8'hFF;
			14'd14068: ff_rdata <= 8'hFF;
			14'd14069: ff_rdata <= 8'hFF;
			14'd14070: ff_rdata <= 8'hFF;
			14'd14071: ff_rdata <= 8'hFF;
			14'd14072: ff_rdata <= 8'hFF;
			14'd14073: ff_rdata <= 8'hFF;
			14'd14074: ff_rdata <= 8'hFF;
			14'd14075: ff_rdata <= 8'hFF;
			14'd14076: ff_rdata <= 8'hFF;
			14'd14077: ff_rdata <= 8'hFF;
			14'd14078: ff_rdata <= 8'hFF;
			14'd14079: ff_rdata <= 8'hFF;
			14'd14080: ff_rdata <= 8'hFF;
			14'd14081: ff_rdata <= 8'hFF;
			14'd14082: ff_rdata <= 8'hFF;
			14'd14083: ff_rdata <= 8'hFF;
			14'd14084: ff_rdata <= 8'hFF;
			14'd14085: ff_rdata <= 8'hFF;
			14'd14086: ff_rdata <= 8'hFF;
			14'd14087: ff_rdata <= 8'hFF;
			14'd14088: ff_rdata <= 8'hFF;
			14'd14089: ff_rdata <= 8'hFF;
			14'd14090: ff_rdata <= 8'hFF;
			14'd14091: ff_rdata <= 8'hFF;
			14'd14092: ff_rdata <= 8'hFF;
			14'd14093: ff_rdata <= 8'hFF;
			14'd14094: ff_rdata <= 8'hFF;
			14'd14095: ff_rdata <= 8'hFF;
			14'd14096: ff_rdata <= 8'hFF;
			14'd14097: ff_rdata <= 8'hFF;
			14'd14098: ff_rdata <= 8'hFF;
			14'd14099: ff_rdata <= 8'hFF;
			14'd14100: ff_rdata <= 8'hFF;
			14'd14101: ff_rdata <= 8'hFF;
			14'd14102: ff_rdata <= 8'hFF;
			14'd14103: ff_rdata <= 8'hFF;
			14'd14104: ff_rdata <= 8'hFF;
			14'd14105: ff_rdata <= 8'hFF;
			14'd14106: ff_rdata <= 8'hFF;
			14'd14107: ff_rdata <= 8'hFF;
			14'd14108: ff_rdata <= 8'hFF;
			14'd14109: ff_rdata <= 8'hFF;
			14'd14110: ff_rdata <= 8'hFF;
			14'd14111: ff_rdata <= 8'hFF;
			14'd14112: ff_rdata <= 8'hFF;
			14'd14113: ff_rdata <= 8'hFF;
			14'd14114: ff_rdata <= 8'hFF;
			14'd14115: ff_rdata <= 8'hFF;
			14'd14116: ff_rdata <= 8'hFF;
			14'd14117: ff_rdata <= 8'hFF;
			14'd14118: ff_rdata <= 8'hFF;
			14'd14119: ff_rdata <= 8'hFF;
			14'd14120: ff_rdata <= 8'hFF;
			14'd14121: ff_rdata <= 8'hFF;
			14'd14122: ff_rdata <= 8'hFF;
			14'd14123: ff_rdata <= 8'hFF;
			14'd14124: ff_rdata <= 8'hFF;
			14'd14125: ff_rdata <= 8'hFF;
			14'd14126: ff_rdata <= 8'hFF;
			14'd14127: ff_rdata <= 8'hFF;
			14'd14128: ff_rdata <= 8'hFF;
			14'd14129: ff_rdata <= 8'hFF;
			14'd14130: ff_rdata <= 8'hFF;
			14'd14131: ff_rdata <= 8'hFF;
			14'd14132: ff_rdata <= 8'hFF;
			14'd14133: ff_rdata <= 8'hFF;
			14'd14134: ff_rdata <= 8'hFF;
			14'd14135: ff_rdata <= 8'hFF;
			14'd14136: ff_rdata <= 8'hFF;
			14'd14137: ff_rdata <= 8'hFF;
			14'd14138: ff_rdata <= 8'hFF;
			14'd14139: ff_rdata <= 8'hFF;
			14'd14140: ff_rdata <= 8'hFF;
			14'd14141: ff_rdata <= 8'hFF;
			14'd14142: ff_rdata <= 8'hFF;
			14'd14143: ff_rdata <= 8'hFF;
			14'd14144: ff_rdata <= 8'hFF;
			14'd14145: ff_rdata <= 8'hFF;
			14'd14146: ff_rdata <= 8'hFF;
			14'd14147: ff_rdata <= 8'hFF;
			14'd14148: ff_rdata <= 8'hFF;
			14'd14149: ff_rdata <= 8'hFF;
			14'd14150: ff_rdata <= 8'hFF;
			14'd14151: ff_rdata <= 8'hFF;
			14'd14152: ff_rdata <= 8'hFF;
			14'd14153: ff_rdata <= 8'hFF;
			14'd14154: ff_rdata <= 8'hFF;
			14'd14155: ff_rdata <= 8'hFF;
			14'd14156: ff_rdata <= 8'hFF;
			14'd14157: ff_rdata <= 8'hFF;
			14'd14158: ff_rdata <= 8'hFF;
			14'd14159: ff_rdata <= 8'hFF;
			14'd14160: ff_rdata <= 8'hFF;
			14'd14161: ff_rdata <= 8'hFF;
			14'd14162: ff_rdata <= 8'hFF;
			14'd14163: ff_rdata <= 8'hFF;
			14'd14164: ff_rdata <= 8'hFF;
			14'd14165: ff_rdata <= 8'hFF;
			14'd14166: ff_rdata <= 8'hFF;
			14'd14167: ff_rdata <= 8'hFF;
			14'd14168: ff_rdata <= 8'hFF;
			14'd14169: ff_rdata <= 8'hFF;
			14'd14170: ff_rdata <= 8'hFF;
			14'd14171: ff_rdata <= 8'hFF;
			14'd14172: ff_rdata <= 8'hFF;
			14'd14173: ff_rdata <= 8'hFF;
			14'd14174: ff_rdata <= 8'hFF;
			14'd14175: ff_rdata <= 8'hFF;
			14'd14176: ff_rdata <= 8'hFF;
			14'd14177: ff_rdata <= 8'hFF;
			14'd14178: ff_rdata <= 8'hFF;
			14'd14179: ff_rdata <= 8'hFF;
			14'd14180: ff_rdata <= 8'hFF;
			14'd14181: ff_rdata <= 8'hFF;
			14'd14182: ff_rdata <= 8'hFF;
			14'd14183: ff_rdata <= 8'hFF;
			14'd14184: ff_rdata <= 8'hFF;
			14'd14185: ff_rdata <= 8'hFF;
			14'd14186: ff_rdata <= 8'hFF;
			14'd14187: ff_rdata <= 8'hFF;
			14'd14188: ff_rdata <= 8'hFF;
			14'd14189: ff_rdata <= 8'hFF;
			14'd14190: ff_rdata <= 8'hFF;
			14'd14191: ff_rdata <= 8'hFF;
			14'd14192: ff_rdata <= 8'hFF;
			14'd14193: ff_rdata <= 8'hFF;
			14'd14194: ff_rdata <= 8'hFF;
			14'd14195: ff_rdata <= 8'hFF;
			14'd14196: ff_rdata <= 8'hFF;
			14'd14197: ff_rdata <= 8'hFF;
			14'd14198: ff_rdata <= 8'hFF;
			14'd14199: ff_rdata <= 8'hFF;
			14'd14200: ff_rdata <= 8'hFF;
			14'd14201: ff_rdata <= 8'hFF;
			14'd14202: ff_rdata <= 8'hFF;
			14'd14203: ff_rdata <= 8'hFF;
			14'd14204: ff_rdata <= 8'hFF;
			14'd14205: ff_rdata <= 8'hFF;
			14'd14206: ff_rdata <= 8'hFF;
			14'd14207: ff_rdata <= 8'hFF;
			14'd14208: ff_rdata <= 8'hFF;
			14'd14209: ff_rdata <= 8'hFF;
			14'd14210: ff_rdata <= 8'hFF;
			14'd14211: ff_rdata <= 8'hFF;
			14'd14212: ff_rdata <= 8'hFF;
			14'd14213: ff_rdata <= 8'hFF;
			14'd14214: ff_rdata <= 8'hFF;
			14'd14215: ff_rdata <= 8'hFF;
			14'd14216: ff_rdata <= 8'hFF;
			14'd14217: ff_rdata <= 8'hFF;
			14'd14218: ff_rdata <= 8'hFF;
			14'd14219: ff_rdata <= 8'hFF;
			14'd14220: ff_rdata <= 8'hFF;
			14'd14221: ff_rdata <= 8'hFF;
			14'd14222: ff_rdata <= 8'hFF;
			14'd14223: ff_rdata <= 8'hFF;
			14'd14224: ff_rdata <= 8'hFF;
			14'd14225: ff_rdata <= 8'hFF;
			14'd14226: ff_rdata <= 8'hFF;
			14'd14227: ff_rdata <= 8'hFF;
			14'd14228: ff_rdata <= 8'hFF;
			14'd14229: ff_rdata <= 8'hFF;
			14'd14230: ff_rdata <= 8'hFF;
			14'd14231: ff_rdata <= 8'hFF;
			14'd14232: ff_rdata <= 8'hFF;
			14'd14233: ff_rdata <= 8'hFF;
			14'd14234: ff_rdata <= 8'hFF;
			14'd14235: ff_rdata <= 8'hFF;
			14'd14236: ff_rdata <= 8'hFF;
			14'd14237: ff_rdata <= 8'hFF;
			14'd14238: ff_rdata <= 8'hFF;
			14'd14239: ff_rdata <= 8'hFF;
			14'd14240: ff_rdata <= 8'hFF;
			14'd14241: ff_rdata <= 8'hFF;
			14'd14242: ff_rdata <= 8'hFF;
			14'd14243: ff_rdata <= 8'hFF;
			14'd14244: ff_rdata <= 8'hFF;
			14'd14245: ff_rdata <= 8'hFF;
			14'd14246: ff_rdata <= 8'hFF;
			14'd14247: ff_rdata <= 8'hFF;
			14'd14248: ff_rdata <= 8'hFF;
			14'd14249: ff_rdata <= 8'hFF;
			14'd14250: ff_rdata <= 8'hFF;
			14'd14251: ff_rdata <= 8'hFF;
			14'd14252: ff_rdata <= 8'hFF;
			14'd14253: ff_rdata <= 8'hFF;
			14'd14254: ff_rdata <= 8'hFF;
			14'd14255: ff_rdata <= 8'hFF;
			14'd14256: ff_rdata <= 8'hFF;
			14'd14257: ff_rdata <= 8'hFF;
			14'd14258: ff_rdata <= 8'hFF;
			14'd14259: ff_rdata <= 8'hFF;
			14'd14260: ff_rdata <= 8'hFF;
			14'd14261: ff_rdata <= 8'hFF;
			14'd14262: ff_rdata <= 8'hFF;
			14'd14263: ff_rdata <= 8'hFF;
			14'd14264: ff_rdata <= 8'hFF;
			14'd14265: ff_rdata <= 8'hFF;
			14'd14266: ff_rdata <= 8'hFF;
			14'd14267: ff_rdata <= 8'hFF;
			14'd14268: ff_rdata <= 8'hFF;
			14'd14269: ff_rdata <= 8'hFF;
			14'd14270: ff_rdata <= 8'hFF;
			14'd14271: ff_rdata <= 8'hFF;
			14'd14272: ff_rdata <= 8'hFF;
			14'd14273: ff_rdata <= 8'hFF;
			14'd14274: ff_rdata <= 8'hFF;
			14'd14275: ff_rdata <= 8'hFF;
			14'd14276: ff_rdata <= 8'hFF;
			14'd14277: ff_rdata <= 8'hFF;
			14'd14278: ff_rdata <= 8'hFF;
			14'd14279: ff_rdata <= 8'hFF;
			14'd14280: ff_rdata <= 8'hFF;
			14'd14281: ff_rdata <= 8'hFF;
			14'd14282: ff_rdata <= 8'hFF;
			14'd14283: ff_rdata <= 8'hFF;
			14'd14284: ff_rdata <= 8'hFF;
			14'd14285: ff_rdata <= 8'hFF;
			14'd14286: ff_rdata <= 8'hFF;
			14'd14287: ff_rdata <= 8'hFF;
			14'd14288: ff_rdata <= 8'hFF;
			14'd14289: ff_rdata <= 8'hFF;
			14'd14290: ff_rdata <= 8'hFF;
			14'd14291: ff_rdata <= 8'hFF;
			14'd14292: ff_rdata <= 8'hFF;
			14'd14293: ff_rdata <= 8'hFF;
			14'd14294: ff_rdata <= 8'hFF;
			14'd14295: ff_rdata <= 8'hFF;
			14'd14296: ff_rdata <= 8'hFF;
			14'd14297: ff_rdata <= 8'hFF;
			14'd14298: ff_rdata <= 8'hFF;
			14'd14299: ff_rdata <= 8'hFF;
			14'd14300: ff_rdata <= 8'hFF;
			14'd14301: ff_rdata <= 8'hFF;
			14'd14302: ff_rdata <= 8'hFF;
			14'd14303: ff_rdata <= 8'hFF;
			14'd14304: ff_rdata <= 8'hFF;
			14'd14305: ff_rdata <= 8'hFF;
			14'd14306: ff_rdata <= 8'hFF;
			14'd14307: ff_rdata <= 8'hFF;
			14'd14308: ff_rdata <= 8'hFF;
			14'd14309: ff_rdata <= 8'hFF;
			14'd14310: ff_rdata <= 8'hFF;
			14'd14311: ff_rdata <= 8'hFF;
			14'd14312: ff_rdata <= 8'hFF;
			14'd14313: ff_rdata <= 8'hFF;
			14'd14314: ff_rdata <= 8'hFF;
			14'd14315: ff_rdata <= 8'hFF;
			14'd14316: ff_rdata <= 8'hFF;
			14'd14317: ff_rdata <= 8'hFF;
			14'd14318: ff_rdata <= 8'hFF;
			14'd14319: ff_rdata <= 8'hFF;
			14'd14320: ff_rdata <= 8'hFF;
			14'd14321: ff_rdata <= 8'hFF;
			14'd14322: ff_rdata <= 8'hFF;
			14'd14323: ff_rdata <= 8'hFF;
			14'd14324: ff_rdata <= 8'hFF;
			14'd14325: ff_rdata <= 8'hFF;
			14'd14326: ff_rdata <= 8'hFF;
			14'd14327: ff_rdata <= 8'hFF;
			14'd14328: ff_rdata <= 8'hFF;
			14'd14329: ff_rdata <= 8'hFF;
			14'd14330: ff_rdata <= 8'hFF;
			14'd14331: ff_rdata <= 8'hFF;
			14'd14332: ff_rdata <= 8'hFF;
			14'd14333: ff_rdata <= 8'hFF;
			14'd14334: ff_rdata <= 8'hFF;
			14'd14335: ff_rdata <= 8'hFF;
			14'd14336: ff_rdata <= 8'hFF;
			14'd14337: ff_rdata <= 8'hFF;
			14'd14338: ff_rdata <= 8'hFF;
			14'd14339: ff_rdata <= 8'hFF;
			14'd14340: ff_rdata <= 8'hFF;
			14'd14341: ff_rdata <= 8'hFF;
			14'd14342: ff_rdata <= 8'hFF;
			14'd14343: ff_rdata <= 8'hFF;
			14'd14344: ff_rdata <= 8'hFF;
			14'd14345: ff_rdata <= 8'hFF;
			14'd14346: ff_rdata <= 8'hFF;
			14'd14347: ff_rdata <= 8'hFF;
			14'd14348: ff_rdata <= 8'hFF;
			14'd14349: ff_rdata <= 8'hFF;
			14'd14350: ff_rdata <= 8'hFF;
			14'd14351: ff_rdata <= 8'hFF;
			14'd14352: ff_rdata <= 8'hFF;
			14'd14353: ff_rdata <= 8'hFF;
			14'd14354: ff_rdata <= 8'hFF;
			14'd14355: ff_rdata <= 8'hFF;
			14'd14356: ff_rdata <= 8'hFF;
			14'd14357: ff_rdata <= 8'hFF;
			14'd14358: ff_rdata <= 8'hFF;
			14'd14359: ff_rdata <= 8'hFF;
			14'd14360: ff_rdata <= 8'hFF;
			14'd14361: ff_rdata <= 8'hFF;
			14'd14362: ff_rdata <= 8'hFF;
			14'd14363: ff_rdata <= 8'hFF;
			14'd14364: ff_rdata <= 8'hFF;
			14'd14365: ff_rdata <= 8'hFF;
			14'd14366: ff_rdata <= 8'hFF;
			14'd14367: ff_rdata <= 8'hFF;
			14'd14368: ff_rdata <= 8'hFF;
			14'd14369: ff_rdata <= 8'hFF;
			14'd14370: ff_rdata <= 8'hFF;
			14'd14371: ff_rdata <= 8'hFF;
			14'd14372: ff_rdata <= 8'hFF;
			14'd14373: ff_rdata <= 8'hFF;
			14'd14374: ff_rdata <= 8'hFF;
			14'd14375: ff_rdata <= 8'hFF;
			14'd14376: ff_rdata <= 8'hFF;
			14'd14377: ff_rdata <= 8'hFF;
			14'd14378: ff_rdata <= 8'hFF;
			14'd14379: ff_rdata <= 8'hFF;
			14'd14380: ff_rdata <= 8'hFF;
			14'd14381: ff_rdata <= 8'hFF;
			14'd14382: ff_rdata <= 8'hFF;
			14'd14383: ff_rdata <= 8'hFF;
			14'd14384: ff_rdata <= 8'hFF;
			14'd14385: ff_rdata <= 8'hFF;
			14'd14386: ff_rdata <= 8'hFF;
			14'd14387: ff_rdata <= 8'hFF;
			14'd14388: ff_rdata <= 8'hFF;
			14'd14389: ff_rdata <= 8'hFF;
			14'd14390: ff_rdata <= 8'hFF;
			14'd14391: ff_rdata <= 8'hFF;
			14'd14392: ff_rdata <= 8'hFF;
			14'd14393: ff_rdata <= 8'hFF;
			14'd14394: ff_rdata <= 8'hFF;
			14'd14395: ff_rdata <= 8'hFF;
			14'd14396: ff_rdata <= 8'hFF;
			14'd14397: ff_rdata <= 8'hFF;
			14'd14398: ff_rdata <= 8'hFF;
			14'd14399: ff_rdata <= 8'hFF;
			14'd14400: ff_rdata <= 8'hFF;
			14'd14401: ff_rdata <= 8'hFF;
			14'd14402: ff_rdata <= 8'hFF;
			14'd14403: ff_rdata <= 8'hFF;
			14'd14404: ff_rdata <= 8'hFF;
			14'd14405: ff_rdata <= 8'hFF;
			14'd14406: ff_rdata <= 8'hFF;
			14'd14407: ff_rdata <= 8'hFF;
			14'd14408: ff_rdata <= 8'hFF;
			14'd14409: ff_rdata <= 8'hFF;
			14'd14410: ff_rdata <= 8'hFF;
			14'd14411: ff_rdata <= 8'hFF;
			14'd14412: ff_rdata <= 8'hFF;
			14'd14413: ff_rdata <= 8'hFF;
			14'd14414: ff_rdata <= 8'hFF;
			14'd14415: ff_rdata <= 8'hFF;
			14'd14416: ff_rdata <= 8'hFF;
			14'd14417: ff_rdata <= 8'hFF;
			14'd14418: ff_rdata <= 8'hFF;
			14'd14419: ff_rdata <= 8'hFF;
			14'd14420: ff_rdata <= 8'hFF;
			14'd14421: ff_rdata <= 8'hFF;
			14'd14422: ff_rdata <= 8'hFF;
			14'd14423: ff_rdata <= 8'hFF;
			14'd14424: ff_rdata <= 8'hFF;
			14'd14425: ff_rdata <= 8'hFF;
			14'd14426: ff_rdata <= 8'hFF;
			14'd14427: ff_rdata <= 8'hFF;
			14'd14428: ff_rdata <= 8'hFF;
			14'd14429: ff_rdata <= 8'hFF;
			14'd14430: ff_rdata <= 8'hFF;
			14'd14431: ff_rdata <= 8'hFF;
			14'd14432: ff_rdata <= 8'hFF;
			14'd14433: ff_rdata <= 8'hFF;
			14'd14434: ff_rdata <= 8'hFF;
			14'd14435: ff_rdata <= 8'hFF;
			14'd14436: ff_rdata <= 8'hFF;
			14'd14437: ff_rdata <= 8'hFF;
			14'd14438: ff_rdata <= 8'hFF;
			14'd14439: ff_rdata <= 8'hFF;
			14'd14440: ff_rdata <= 8'hFF;
			14'd14441: ff_rdata <= 8'hFF;
			14'd14442: ff_rdata <= 8'hFF;
			14'd14443: ff_rdata <= 8'hFF;
			14'd14444: ff_rdata <= 8'hFF;
			14'd14445: ff_rdata <= 8'hFF;
			14'd14446: ff_rdata <= 8'hFF;
			14'd14447: ff_rdata <= 8'hFF;
			14'd14448: ff_rdata <= 8'hFF;
			14'd14449: ff_rdata <= 8'hFF;
			14'd14450: ff_rdata <= 8'hFF;
			14'd14451: ff_rdata <= 8'hFF;
			14'd14452: ff_rdata <= 8'hFF;
			14'd14453: ff_rdata <= 8'hFF;
			14'd14454: ff_rdata <= 8'hFF;
			14'd14455: ff_rdata <= 8'hFF;
			14'd14456: ff_rdata <= 8'hFF;
			14'd14457: ff_rdata <= 8'hFF;
			14'd14458: ff_rdata <= 8'hFF;
			14'd14459: ff_rdata <= 8'hFF;
			14'd14460: ff_rdata <= 8'hFF;
			14'd14461: ff_rdata <= 8'hFF;
			14'd14462: ff_rdata <= 8'hFF;
			14'd14463: ff_rdata <= 8'hFF;
			14'd14464: ff_rdata <= 8'hFF;
			14'd14465: ff_rdata <= 8'hFF;
			14'd14466: ff_rdata <= 8'hFF;
			14'd14467: ff_rdata <= 8'hFF;
			14'd14468: ff_rdata <= 8'hFF;
			14'd14469: ff_rdata <= 8'hFF;
			14'd14470: ff_rdata <= 8'hFF;
			14'd14471: ff_rdata <= 8'hFF;
			14'd14472: ff_rdata <= 8'hFF;
			14'd14473: ff_rdata <= 8'hFF;
			14'd14474: ff_rdata <= 8'hFF;
			14'd14475: ff_rdata <= 8'hFF;
			14'd14476: ff_rdata <= 8'hFF;
			14'd14477: ff_rdata <= 8'hFF;
			14'd14478: ff_rdata <= 8'hFF;
			14'd14479: ff_rdata <= 8'hFF;
			14'd14480: ff_rdata <= 8'hFF;
			14'd14481: ff_rdata <= 8'hFF;
			14'd14482: ff_rdata <= 8'hFF;
			14'd14483: ff_rdata <= 8'hFF;
			14'd14484: ff_rdata <= 8'hFF;
			14'd14485: ff_rdata <= 8'hFF;
			14'd14486: ff_rdata <= 8'hFF;
			14'd14487: ff_rdata <= 8'hFF;
			14'd14488: ff_rdata <= 8'hFF;
			14'd14489: ff_rdata <= 8'hFF;
			14'd14490: ff_rdata <= 8'hFF;
			14'd14491: ff_rdata <= 8'hFF;
			14'd14492: ff_rdata <= 8'hFF;
			14'd14493: ff_rdata <= 8'hFF;
			14'd14494: ff_rdata <= 8'hFF;
			14'd14495: ff_rdata <= 8'hFF;
			14'd14496: ff_rdata <= 8'hFF;
			14'd14497: ff_rdata <= 8'hFF;
			14'd14498: ff_rdata <= 8'hFF;
			14'd14499: ff_rdata <= 8'hFF;
			14'd14500: ff_rdata <= 8'hFF;
			14'd14501: ff_rdata <= 8'hFF;
			14'd14502: ff_rdata <= 8'hFF;
			14'd14503: ff_rdata <= 8'hFF;
			14'd14504: ff_rdata <= 8'hFF;
			14'd14505: ff_rdata <= 8'hFF;
			14'd14506: ff_rdata <= 8'hFF;
			14'd14507: ff_rdata <= 8'hFF;
			14'd14508: ff_rdata <= 8'hFF;
			14'd14509: ff_rdata <= 8'hFF;
			14'd14510: ff_rdata <= 8'hFF;
			14'd14511: ff_rdata <= 8'hFF;
			14'd14512: ff_rdata <= 8'hFF;
			14'd14513: ff_rdata <= 8'hFF;
			14'd14514: ff_rdata <= 8'hFF;
			14'd14515: ff_rdata <= 8'hFF;
			14'd14516: ff_rdata <= 8'hFF;
			14'd14517: ff_rdata <= 8'hFF;
			14'd14518: ff_rdata <= 8'hFF;
			14'd14519: ff_rdata <= 8'hFF;
			14'd14520: ff_rdata <= 8'hFF;
			14'd14521: ff_rdata <= 8'hFF;
			14'd14522: ff_rdata <= 8'hFF;
			14'd14523: ff_rdata <= 8'hFF;
			14'd14524: ff_rdata <= 8'hFF;
			14'd14525: ff_rdata <= 8'hFF;
			14'd14526: ff_rdata <= 8'hFF;
			14'd14527: ff_rdata <= 8'hFF;
			14'd14528: ff_rdata <= 8'hFF;
			14'd14529: ff_rdata <= 8'hFF;
			14'd14530: ff_rdata <= 8'hFF;
			14'd14531: ff_rdata <= 8'hFF;
			14'd14532: ff_rdata <= 8'hFF;
			14'd14533: ff_rdata <= 8'hFF;
			14'd14534: ff_rdata <= 8'hFF;
			14'd14535: ff_rdata <= 8'hFF;
			14'd14536: ff_rdata <= 8'hFF;
			14'd14537: ff_rdata <= 8'hFF;
			14'd14538: ff_rdata <= 8'hFF;
			14'd14539: ff_rdata <= 8'hFF;
			14'd14540: ff_rdata <= 8'hFF;
			14'd14541: ff_rdata <= 8'hFF;
			14'd14542: ff_rdata <= 8'hFF;
			14'd14543: ff_rdata <= 8'hFF;
			14'd14544: ff_rdata <= 8'hFF;
			14'd14545: ff_rdata <= 8'hFF;
			14'd14546: ff_rdata <= 8'hFF;
			14'd14547: ff_rdata <= 8'hFF;
			14'd14548: ff_rdata <= 8'hFF;
			14'd14549: ff_rdata <= 8'hFF;
			14'd14550: ff_rdata <= 8'hFF;
			14'd14551: ff_rdata <= 8'hFF;
			14'd14552: ff_rdata <= 8'hFF;
			14'd14553: ff_rdata <= 8'hFF;
			14'd14554: ff_rdata <= 8'hFF;
			14'd14555: ff_rdata <= 8'hFF;
			14'd14556: ff_rdata <= 8'hFF;
			14'd14557: ff_rdata <= 8'hFF;
			14'd14558: ff_rdata <= 8'hFF;
			14'd14559: ff_rdata <= 8'hFF;
			14'd14560: ff_rdata <= 8'hFF;
			14'd14561: ff_rdata <= 8'hFF;
			14'd14562: ff_rdata <= 8'hFF;
			14'd14563: ff_rdata <= 8'hFF;
			14'd14564: ff_rdata <= 8'hFF;
			14'd14565: ff_rdata <= 8'hFF;
			14'd14566: ff_rdata <= 8'hFF;
			14'd14567: ff_rdata <= 8'hFF;
			14'd14568: ff_rdata <= 8'hFF;
			14'd14569: ff_rdata <= 8'hFF;
			14'd14570: ff_rdata <= 8'hFF;
			14'd14571: ff_rdata <= 8'hFF;
			14'd14572: ff_rdata <= 8'hFF;
			14'd14573: ff_rdata <= 8'hFF;
			14'd14574: ff_rdata <= 8'hFF;
			14'd14575: ff_rdata <= 8'hFF;
			14'd14576: ff_rdata <= 8'hFF;
			14'd14577: ff_rdata <= 8'hFF;
			14'd14578: ff_rdata <= 8'hFF;
			14'd14579: ff_rdata <= 8'hFF;
			14'd14580: ff_rdata <= 8'hFF;
			14'd14581: ff_rdata <= 8'hFF;
			14'd14582: ff_rdata <= 8'hFF;
			14'd14583: ff_rdata <= 8'hFF;
			14'd14584: ff_rdata <= 8'hFF;
			14'd14585: ff_rdata <= 8'hFF;
			14'd14586: ff_rdata <= 8'hFF;
			14'd14587: ff_rdata <= 8'hFF;
			14'd14588: ff_rdata <= 8'hFF;
			14'd14589: ff_rdata <= 8'hFF;
			14'd14590: ff_rdata <= 8'hFF;
			14'd14591: ff_rdata <= 8'hFF;
			14'd14592: ff_rdata <= 8'hFF;
			14'd14593: ff_rdata <= 8'hFF;
			14'd14594: ff_rdata <= 8'hFF;
			14'd14595: ff_rdata <= 8'hFF;
			14'd14596: ff_rdata <= 8'hFF;
			14'd14597: ff_rdata <= 8'hFF;
			14'd14598: ff_rdata <= 8'hFF;
			14'd14599: ff_rdata <= 8'hFF;
			14'd14600: ff_rdata <= 8'hFF;
			14'd14601: ff_rdata <= 8'hFF;
			14'd14602: ff_rdata <= 8'hFF;
			14'd14603: ff_rdata <= 8'hFF;
			14'd14604: ff_rdata <= 8'hFF;
			14'd14605: ff_rdata <= 8'hFF;
			14'd14606: ff_rdata <= 8'hFF;
			14'd14607: ff_rdata <= 8'hFF;
			14'd14608: ff_rdata <= 8'hFF;
			14'd14609: ff_rdata <= 8'hFF;
			14'd14610: ff_rdata <= 8'hFF;
			14'd14611: ff_rdata <= 8'hFF;
			14'd14612: ff_rdata <= 8'hFF;
			14'd14613: ff_rdata <= 8'hFF;
			14'd14614: ff_rdata <= 8'hFF;
			14'd14615: ff_rdata <= 8'hFF;
			14'd14616: ff_rdata <= 8'hFF;
			14'd14617: ff_rdata <= 8'hFF;
			14'd14618: ff_rdata <= 8'hFF;
			14'd14619: ff_rdata <= 8'hFF;
			14'd14620: ff_rdata <= 8'hFF;
			14'd14621: ff_rdata <= 8'hFF;
			14'd14622: ff_rdata <= 8'hFF;
			14'd14623: ff_rdata <= 8'hFF;
			14'd14624: ff_rdata <= 8'hFF;
			14'd14625: ff_rdata <= 8'hFF;
			14'd14626: ff_rdata <= 8'hFF;
			14'd14627: ff_rdata <= 8'hFF;
			14'd14628: ff_rdata <= 8'hFF;
			14'd14629: ff_rdata <= 8'hFF;
			14'd14630: ff_rdata <= 8'hFF;
			14'd14631: ff_rdata <= 8'hFF;
			14'd14632: ff_rdata <= 8'hFF;
			14'd14633: ff_rdata <= 8'hFF;
			14'd14634: ff_rdata <= 8'hFF;
			14'd14635: ff_rdata <= 8'hFF;
			14'd14636: ff_rdata <= 8'hFF;
			14'd14637: ff_rdata <= 8'hFF;
			14'd14638: ff_rdata <= 8'hFF;
			14'd14639: ff_rdata <= 8'hFF;
			14'd14640: ff_rdata <= 8'hFF;
			14'd14641: ff_rdata <= 8'hFF;
			14'd14642: ff_rdata <= 8'hFF;
			14'd14643: ff_rdata <= 8'hFF;
			14'd14644: ff_rdata <= 8'hFF;
			14'd14645: ff_rdata <= 8'hFF;
			14'd14646: ff_rdata <= 8'hFF;
			14'd14647: ff_rdata <= 8'hFF;
			14'd14648: ff_rdata <= 8'hFF;
			14'd14649: ff_rdata <= 8'hFF;
			14'd14650: ff_rdata <= 8'hFF;
			14'd14651: ff_rdata <= 8'hFF;
			14'd14652: ff_rdata <= 8'hFF;
			14'd14653: ff_rdata <= 8'hFF;
			14'd14654: ff_rdata <= 8'hFF;
			14'd14655: ff_rdata <= 8'hFF;
			14'd14656: ff_rdata <= 8'hFF;
			14'd14657: ff_rdata <= 8'hFF;
			14'd14658: ff_rdata <= 8'hFF;
			14'd14659: ff_rdata <= 8'hFF;
			14'd14660: ff_rdata <= 8'hFF;
			14'd14661: ff_rdata <= 8'hFF;
			14'd14662: ff_rdata <= 8'hFF;
			14'd14663: ff_rdata <= 8'hFF;
			14'd14664: ff_rdata <= 8'hFF;
			14'd14665: ff_rdata <= 8'hFF;
			14'd14666: ff_rdata <= 8'hFF;
			14'd14667: ff_rdata <= 8'hFF;
			14'd14668: ff_rdata <= 8'hFF;
			14'd14669: ff_rdata <= 8'hFF;
			14'd14670: ff_rdata <= 8'hFF;
			14'd14671: ff_rdata <= 8'hFF;
			14'd14672: ff_rdata <= 8'hFF;
			14'd14673: ff_rdata <= 8'hFF;
			14'd14674: ff_rdata <= 8'hFF;
			14'd14675: ff_rdata <= 8'hFF;
			14'd14676: ff_rdata <= 8'hFF;
			14'd14677: ff_rdata <= 8'hFF;
			14'd14678: ff_rdata <= 8'hFF;
			14'd14679: ff_rdata <= 8'hFF;
			14'd14680: ff_rdata <= 8'hFF;
			14'd14681: ff_rdata <= 8'hFF;
			14'd14682: ff_rdata <= 8'hFF;
			14'd14683: ff_rdata <= 8'hFF;
			14'd14684: ff_rdata <= 8'hFF;
			14'd14685: ff_rdata <= 8'hFF;
			14'd14686: ff_rdata <= 8'hFF;
			14'd14687: ff_rdata <= 8'hFF;
			14'd14688: ff_rdata <= 8'hFF;
			14'd14689: ff_rdata <= 8'hFF;
			14'd14690: ff_rdata <= 8'hFF;
			14'd14691: ff_rdata <= 8'hFF;
			14'd14692: ff_rdata <= 8'hFF;
			14'd14693: ff_rdata <= 8'hFF;
			14'd14694: ff_rdata <= 8'hFF;
			14'd14695: ff_rdata <= 8'hFF;
			14'd14696: ff_rdata <= 8'hFF;
			14'd14697: ff_rdata <= 8'hFF;
			14'd14698: ff_rdata <= 8'hFF;
			14'd14699: ff_rdata <= 8'hFF;
			14'd14700: ff_rdata <= 8'hFF;
			14'd14701: ff_rdata <= 8'hFF;
			14'd14702: ff_rdata <= 8'hFF;
			14'd14703: ff_rdata <= 8'hFF;
			14'd14704: ff_rdata <= 8'hFF;
			14'd14705: ff_rdata <= 8'hFF;
			14'd14706: ff_rdata <= 8'hFF;
			14'd14707: ff_rdata <= 8'hFF;
			14'd14708: ff_rdata <= 8'hFF;
			14'd14709: ff_rdata <= 8'hFF;
			14'd14710: ff_rdata <= 8'hFF;
			14'd14711: ff_rdata <= 8'hFF;
			14'd14712: ff_rdata <= 8'hFF;
			14'd14713: ff_rdata <= 8'hFF;
			14'd14714: ff_rdata <= 8'hFF;
			14'd14715: ff_rdata <= 8'hFF;
			14'd14716: ff_rdata <= 8'hFF;
			14'd14717: ff_rdata <= 8'hFF;
			14'd14718: ff_rdata <= 8'hFF;
			14'd14719: ff_rdata <= 8'hFF;
			14'd14720: ff_rdata <= 8'hFF;
			14'd14721: ff_rdata <= 8'hFF;
			14'd14722: ff_rdata <= 8'hFF;
			14'd14723: ff_rdata <= 8'hFF;
			14'd14724: ff_rdata <= 8'hFF;
			14'd14725: ff_rdata <= 8'hFF;
			14'd14726: ff_rdata <= 8'hFF;
			14'd14727: ff_rdata <= 8'hFF;
			14'd14728: ff_rdata <= 8'hFF;
			14'd14729: ff_rdata <= 8'hFF;
			14'd14730: ff_rdata <= 8'hFF;
			14'd14731: ff_rdata <= 8'hFF;
			14'd14732: ff_rdata <= 8'hFF;
			14'd14733: ff_rdata <= 8'hFF;
			14'd14734: ff_rdata <= 8'hFF;
			14'd14735: ff_rdata <= 8'hFF;
			14'd14736: ff_rdata <= 8'hFF;
			14'd14737: ff_rdata <= 8'hFF;
			14'd14738: ff_rdata <= 8'hFF;
			14'd14739: ff_rdata <= 8'hFF;
			14'd14740: ff_rdata <= 8'hFF;
			14'd14741: ff_rdata <= 8'hFF;
			14'd14742: ff_rdata <= 8'hFF;
			14'd14743: ff_rdata <= 8'hFF;
			14'd14744: ff_rdata <= 8'hFF;
			14'd14745: ff_rdata <= 8'hFF;
			14'd14746: ff_rdata <= 8'hFF;
			14'd14747: ff_rdata <= 8'hFF;
			14'd14748: ff_rdata <= 8'hFF;
			14'd14749: ff_rdata <= 8'hFF;
			14'd14750: ff_rdata <= 8'hFF;
			14'd14751: ff_rdata <= 8'hFF;
			14'd14752: ff_rdata <= 8'hFF;
			14'd14753: ff_rdata <= 8'hFF;
			14'd14754: ff_rdata <= 8'hFF;
			14'd14755: ff_rdata <= 8'hFF;
			14'd14756: ff_rdata <= 8'hFF;
			14'd14757: ff_rdata <= 8'hFF;
			14'd14758: ff_rdata <= 8'hFF;
			14'd14759: ff_rdata <= 8'hFF;
			14'd14760: ff_rdata <= 8'hFF;
			14'd14761: ff_rdata <= 8'hFF;
			14'd14762: ff_rdata <= 8'hFF;
			14'd14763: ff_rdata <= 8'hFF;
			14'd14764: ff_rdata <= 8'hFF;
			14'd14765: ff_rdata <= 8'hFF;
			14'd14766: ff_rdata <= 8'hFF;
			14'd14767: ff_rdata <= 8'hFF;
			14'd14768: ff_rdata <= 8'hFF;
			14'd14769: ff_rdata <= 8'hFF;
			14'd14770: ff_rdata <= 8'hFF;
			14'd14771: ff_rdata <= 8'hFF;
			14'd14772: ff_rdata <= 8'hFF;
			14'd14773: ff_rdata <= 8'hFF;
			14'd14774: ff_rdata <= 8'hFF;
			14'd14775: ff_rdata <= 8'hFF;
			14'd14776: ff_rdata <= 8'hFF;
			14'd14777: ff_rdata <= 8'hFF;
			14'd14778: ff_rdata <= 8'hFF;
			14'd14779: ff_rdata <= 8'hFF;
			14'd14780: ff_rdata <= 8'hFF;
			14'd14781: ff_rdata <= 8'hFF;
			14'd14782: ff_rdata <= 8'hFF;
			14'd14783: ff_rdata <= 8'hFF;
			14'd14784: ff_rdata <= 8'hFF;
			14'd14785: ff_rdata <= 8'hFF;
			14'd14786: ff_rdata <= 8'hFF;
			14'd14787: ff_rdata <= 8'hFF;
			14'd14788: ff_rdata <= 8'hFF;
			14'd14789: ff_rdata <= 8'hFF;
			14'd14790: ff_rdata <= 8'hFF;
			14'd14791: ff_rdata <= 8'hFF;
			14'd14792: ff_rdata <= 8'hFF;
			14'd14793: ff_rdata <= 8'hFF;
			14'd14794: ff_rdata <= 8'hFF;
			14'd14795: ff_rdata <= 8'hFF;
			14'd14796: ff_rdata <= 8'hFF;
			14'd14797: ff_rdata <= 8'hFF;
			14'd14798: ff_rdata <= 8'hFF;
			14'd14799: ff_rdata <= 8'hFF;
			14'd14800: ff_rdata <= 8'hFF;
			14'd14801: ff_rdata <= 8'hFF;
			14'd14802: ff_rdata <= 8'hFF;
			14'd14803: ff_rdata <= 8'hFF;
			14'd14804: ff_rdata <= 8'hFF;
			14'd14805: ff_rdata <= 8'hFF;
			14'd14806: ff_rdata <= 8'hFF;
			14'd14807: ff_rdata <= 8'hFF;
			14'd14808: ff_rdata <= 8'hFF;
			14'd14809: ff_rdata <= 8'hFF;
			14'd14810: ff_rdata <= 8'hFF;
			14'd14811: ff_rdata <= 8'hFF;
			14'd14812: ff_rdata <= 8'hFF;
			14'd14813: ff_rdata <= 8'hFF;
			14'd14814: ff_rdata <= 8'hFF;
			14'd14815: ff_rdata <= 8'hFF;
			14'd14816: ff_rdata <= 8'hFF;
			14'd14817: ff_rdata <= 8'hFF;
			14'd14818: ff_rdata <= 8'hFF;
			14'd14819: ff_rdata <= 8'hFF;
			14'd14820: ff_rdata <= 8'hFF;
			14'd14821: ff_rdata <= 8'hFF;
			14'd14822: ff_rdata <= 8'hFF;
			14'd14823: ff_rdata <= 8'hFF;
			14'd14824: ff_rdata <= 8'hFF;
			14'd14825: ff_rdata <= 8'hFF;
			14'd14826: ff_rdata <= 8'hFF;
			14'd14827: ff_rdata <= 8'hFF;
			14'd14828: ff_rdata <= 8'hFF;
			14'd14829: ff_rdata <= 8'hFF;
			14'd14830: ff_rdata <= 8'hFF;
			14'd14831: ff_rdata <= 8'hFF;
			14'd14832: ff_rdata <= 8'hFF;
			14'd14833: ff_rdata <= 8'hFF;
			14'd14834: ff_rdata <= 8'hFF;
			14'd14835: ff_rdata <= 8'hFF;
			14'd14836: ff_rdata <= 8'hFF;
			14'd14837: ff_rdata <= 8'hFF;
			14'd14838: ff_rdata <= 8'hFF;
			14'd14839: ff_rdata <= 8'hFF;
			14'd14840: ff_rdata <= 8'hFF;
			14'd14841: ff_rdata <= 8'hFF;
			14'd14842: ff_rdata <= 8'hFF;
			14'd14843: ff_rdata <= 8'hFF;
			14'd14844: ff_rdata <= 8'hFF;
			14'd14845: ff_rdata <= 8'hFF;
			14'd14846: ff_rdata <= 8'hFF;
			14'd14847: ff_rdata <= 8'hFF;
			14'd14848: ff_rdata <= 8'hFF;
			14'd14849: ff_rdata <= 8'hFF;
			14'd14850: ff_rdata <= 8'hFF;
			14'd14851: ff_rdata <= 8'hFF;
			14'd14852: ff_rdata <= 8'hFF;
			14'd14853: ff_rdata <= 8'hFF;
			14'd14854: ff_rdata <= 8'hFF;
			14'd14855: ff_rdata <= 8'hFF;
			14'd14856: ff_rdata <= 8'hFF;
			14'd14857: ff_rdata <= 8'hFF;
			14'd14858: ff_rdata <= 8'hFF;
			14'd14859: ff_rdata <= 8'hFF;
			14'd14860: ff_rdata <= 8'hFF;
			14'd14861: ff_rdata <= 8'hFF;
			14'd14862: ff_rdata <= 8'hFF;
			14'd14863: ff_rdata <= 8'hFF;
			14'd14864: ff_rdata <= 8'hFF;
			14'd14865: ff_rdata <= 8'hFF;
			14'd14866: ff_rdata <= 8'hFF;
			14'd14867: ff_rdata <= 8'hFF;
			14'd14868: ff_rdata <= 8'hFF;
			14'd14869: ff_rdata <= 8'hFF;
			14'd14870: ff_rdata <= 8'hFF;
			14'd14871: ff_rdata <= 8'hFF;
			14'd14872: ff_rdata <= 8'hFF;
			14'd14873: ff_rdata <= 8'hFF;
			14'd14874: ff_rdata <= 8'hFF;
			14'd14875: ff_rdata <= 8'hFF;
			14'd14876: ff_rdata <= 8'hFF;
			14'd14877: ff_rdata <= 8'hFF;
			14'd14878: ff_rdata <= 8'hFF;
			14'd14879: ff_rdata <= 8'hFF;
			14'd14880: ff_rdata <= 8'hFF;
			14'd14881: ff_rdata <= 8'hFF;
			14'd14882: ff_rdata <= 8'hFF;
			14'd14883: ff_rdata <= 8'hFF;
			14'd14884: ff_rdata <= 8'hFF;
			14'd14885: ff_rdata <= 8'hFF;
			14'd14886: ff_rdata <= 8'hFF;
			14'd14887: ff_rdata <= 8'hFF;
			14'd14888: ff_rdata <= 8'hFF;
			14'd14889: ff_rdata <= 8'hFF;
			14'd14890: ff_rdata <= 8'hFF;
			14'd14891: ff_rdata <= 8'hFF;
			14'd14892: ff_rdata <= 8'hFF;
			14'd14893: ff_rdata <= 8'hFF;
			14'd14894: ff_rdata <= 8'hFF;
			14'd14895: ff_rdata <= 8'hFF;
			14'd14896: ff_rdata <= 8'hFF;
			14'd14897: ff_rdata <= 8'hFF;
			14'd14898: ff_rdata <= 8'hFF;
			14'd14899: ff_rdata <= 8'hFF;
			14'd14900: ff_rdata <= 8'hFF;
			14'd14901: ff_rdata <= 8'hFF;
			14'd14902: ff_rdata <= 8'hFF;
			14'd14903: ff_rdata <= 8'hFF;
			14'd14904: ff_rdata <= 8'hFF;
			14'd14905: ff_rdata <= 8'hFF;
			14'd14906: ff_rdata <= 8'hFF;
			14'd14907: ff_rdata <= 8'hFF;
			14'd14908: ff_rdata <= 8'hFF;
			14'd14909: ff_rdata <= 8'hFF;
			14'd14910: ff_rdata <= 8'hFF;
			14'd14911: ff_rdata <= 8'hFF;
			14'd14912: ff_rdata <= 8'hFF;
			14'd14913: ff_rdata <= 8'hFF;
			14'd14914: ff_rdata <= 8'hFF;
			14'd14915: ff_rdata <= 8'hFF;
			14'd14916: ff_rdata <= 8'hFF;
			14'd14917: ff_rdata <= 8'hFF;
			14'd14918: ff_rdata <= 8'hFF;
			14'd14919: ff_rdata <= 8'hFF;
			14'd14920: ff_rdata <= 8'hFF;
			14'd14921: ff_rdata <= 8'hFF;
			14'd14922: ff_rdata <= 8'hFF;
			14'd14923: ff_rdata <= 8'hFF;
			14'd14924: ff_rdata <= 8'hFF;
			14'd14925: ff_rdata <= 8'hFF;
			14'd14926: ff_rdata <= 8'hFF;
			14'd14927: ff_rdata <= 8'hFF;
			14'd14928: ff_rdata <= 8'hFF;
			14'd14929: ff_rdata <= 8'hFF;
			14'd14930: ff_rdata <= 8'hFF;
			14'd14931: ff_rdata <= 8'hFF;
			14'd14932: ff_rdata <= 8'hFF;
			14'd14933: ff_rdata <= 8'hFF;
			14'd14934: ff_rdata <= 8'hFF;
			14'd14935: ff_rdata <= 8'hFF;
			14'd14936: ff_rdata <= 8'hFF;
			14'd14937: ff_rdata <= 8'hFF;
			14'd14938: ff_rdata <= 8'hFF;
			14'd14939: ff_rdata <= 8'hFF;
			14'd14940: ff_rdata <= 8'hFF;
			14'd14941: ff_rdata <= 8'hFF;
			14'd14942: ff_rdata <= 8'hFF;
			14'd14943: ff_rdata <= 8'hFF;
			14'd14944: ff_rdata <= 8'hFF;
			14'd14945: ff_rdata <= 8'hFF;
			14'd14946: ff_rdata <= 8'hFF;
			14'd14947: ff_rdata <= 8'hFF;
			14'd14948: ff_rdata <= 8'hFF;
			14'd14949: ff_rdata <= 8'hFF;
			14'd14950: ff_rdata <= 8'hFF;
			14'd14951: ff_rdata <= 8'hFF;
			14'd14952: ff_rdata <= 8'hFF;
			14'd14953: ff_rdata <= 8'hFF;
			14'd14954: ff_rdata <= 8'hFF;
			14'd14955: ff_rdata <= 8'hFF;
			14'd14956: ff_rdata <= 8'hFF;
			14'd14957: ff_rdata <= 8'hFF;
			14'd14958: ff_rdata <= 8'hFF;
			14'd14959: ff_rdata <= 8'hFF;
			14'd14960: ff_rdata <= 8'hFF;
			14'd14961: ff_rdata <= 8'hFF;
			14'd14962: ff_rdata <= 8'hFF;
			14'd14963: ff_rdata <= 8'hFF;
			14'd14964: ff_rdata <= 8'hFF;
			14'd14965: ff_rdata <= 8'hFF;
			14'd14966: ff_rdata <= 8'hFF;
			14'd14967: ff_rdata <= 8'hFF;
			14'd14968: ff_rdata <= 8'hFF;
			14'd14969: ff_rdata <= 8'hFF;
			14'd14970: ff_rdata <= 8'hFF;
			14'd14971: ff_rdata <= 8'hFF;
			14'd14972: ff_rdata <= 8'hFF;
			14'd14973: ff_rdata <= 8'hFF;
			14'd14974: ff_rdata <= 8'hFF;
			14'd14975: ff_rdata <= 8'hFF;
			14'd14976: ff_rdata <= 8'hFF;
			14'd14977: ff_rdata <= 8'hFF;
			14'd14978: ff_rdata <= 8'hFF;
			14'd14979: ff_rdata <= 8'hFF;
			14'd14980: ff_rdata <= 8'hFF;
			14'd14981: ff_rdata <= 8'hFF;
			14'd14982: ff_rdata <= 8'hFF;
			14'd14983: ff_rdata <= 8'hFF;
			14'd14984: ff_rdata <= 8'hFF;
			14'd14985: ff_rdata <= 8'hFF;
			14'd14986: ff_rdata <= 8'hFF;
			14'd14987: ff_rdata <= 8'hFF;
			14'd14988: ff_rdata <= 8'hFF;
			14'd14989: ff_rdata <= 8'hFF;
			14'd14990: ff_rdata <= 8'hFF;
			14'd14991: ff_rdata <= 8'hFF;
			14'd14992: ff_rdata <= 8'hFF;
			14'd14993: ff_rdata <= 8'hFF;
			14'd14994: ff_rdata <= 8'hFF;
			14'd14995: ff_rdata <= 8'hFF;
			14'd14996: ff_rdata <= 8'hFF;
			14'd14997: ff_rdata <= 8'hFF;
			14'd14998: ff_rdata <= 8'hFF;
			14'd14999: ff_rdata <= 8'hFF;
			14'd15000: ff_rdata <= 8'hFF;
			14'd15001: ff_rdata <= 8'hFF;
			14'd15002: ff_rdata <= 8'hFF;
			14'd15003: ff_rdata <= 8'hFF;
			14'd15004: ff_rdata <= 8'hFF;
			14'd15005: ff_rdata <= 8'hFF;
			14'd15006: ff_rdata <= 8'hFF;
			14'd15007: ff_rdata <= 8'hFF;
			14'd15008: ff_rdata <= 8'hFF;
			14'd15009: ff_rdata <= 8'hFF;
			14'd15010: ff_rdata <= 8'hFF;
			14'd15011: ff_rdata <= 8'hFF;
			14'd15012: ff_rdata <= 8'hFF;
			14'd15013: ff_rdata <= 8'hFF;
			14'd15014: ff_rdata <= 8'hFF;
			14'd15015: ff_rdata <= 8'hFF;
			14'd15016: ff_rdata <= 8'hFF;
			14'd15017: ff_rdata <= 8'hFF;
			14'd15018: ff_rdata <= 8'hFF;
			14'd15019: ff_rdata <= 8'hFF;
			14'd15020: ff_rdata <= 8'hFF;
			14'd15021: ff_rdata <= 8'hFF;
			14'd15022: ff_rdata <= 8'hFF;
			14'd15023: ff_rdata <= 8'hFF;
			14'd15024: ff_rdata <= 8'hFF;
			14'd15025: ff_rdata <= 8'hFF;
			14'd15026: ff_rdata <= 8'hFF;
			14'd15027: ff_rdata <= 8'hFF;
			14'd15028: ff_rdata <= 8'hFF;
			14'd15029: ff_rdata <= 8'hFF;
			14'd15030: ff_rdata <= 8'hFF;
			14'd15031: ff_rdata <= 8'hFF;
			14'd15032: ff_rdata <= 8'hFF;
			14'd15033: ff_rdata <= 8'hFF;
			14'd15034: ff_rdata <= 8'hFF;
			14'd15035: ff_rdata <= 8'hFF;
			14'd15036: ff_rdata <= 8'hFF;
			14'd15037: ff_rdata <= 8'hFF;
			14'd15038: ff_rdata <= 8'hFF;
			14'd15039: ff_rdata <= 8'hFF;
			14'd15040: ff_rdata <= 8'hFF;
			14'd15041: ff_rdata <= 8'hFF;
			14'd15042: ff_rdata <= 8'hFF;
			14'd15043: ff_rdata <= 8'hFF;
			14'd15044: ff_rdata <= 8'hFF;
			14'd15045: ff_rdata <= 8'hFF;
			14'd15046: ff_rdata <= 8'hFF;
			14'd15047: ff_rdata <= 8'hFF;
			14'd15048: ff_rdata <= 8'hFF;
			14'd15049: ff_rdata <= 8'hFF;
			14'd15050: ff_rdata <= 8'hFF;
			14'd15051: ff_rdata <= 8'hFF;
			14'd15052: ff_rdata <= 8'hFF;
			14'd15053: ff_rdata <= 8'hFF;
			14'd15054: ff_rdata <= 8'hFF;
			14'd15055: ff_rdata <= 8'hFF;
			14'd15056: ff_rdata <= 8'hFF;
			14'd15057: ff_rdata <= 8'hFF;
			14'd15058: ff_rdata <= 8'hFF;
			14'd15059: ff_rdata <= 8'hFF;
			14'd15060: ff_rdata <= 8'hFF;
			14'd15061: ff_rdata <= 8'hFF;
			14'd15062: ff_rdata <= 8'hFF;
			14'd15063: ff_rdata <= 8'hFF;
			14'd15064: ff_rdata <= 8'hFF;
			14'd15065: ff_rdata <= 8'hFF;
			14'd15066: ff_rdata <= 8'hFF;
			14'd15067: ff_rdata <= 8'hFF;
			14'd15068: ff_rdata <= 8'hFF;
			14'd15069: ff_rdata <= 8'hFF;
			14'd15070: ff_rdata <= 8'hFF;
			14'd15071: ff_rdata <= 8'hFF;
			14'd15072: ff_rdata <= 8'hFF;
			14'd15073: ff_rdata <= 8'hFF;
			14'd15074: ff_rdata <= 8'hFF;
			14'd15075: ff_rdata <= 8'hFF;
			14'd15076: ff_rdata <= 8'hFF;
			14'd15077: ff_rdata <= 8'hFF;
			14'd15078: ff_rdata <= 8'hFF;
			14'd15079: ff_rdata <= 8'hFF;
			14'd15080: ff_rdata <= 8'hFF;
			14'd15081: ff_rdata <= 8'hFF;
			14'd15082: ff_rdata <= 8'hFF;
			14'd15083: ff_rdata <= 8'hFF;
			14'd15084: ff_rdata <= 8'hFF;
			14'd15085: ff_rdata <= 8'hFF;
			14'd15086: ff_rdata <= 8'hFF;
			14'd15087: ff_rdata <= 8'hFF;
			14'd15088: ff_rdata <= 8'hFF;
			14'd15089: ff_rdata <= 8'hFF;
			14'd15090: ff_rdata <= 8'hFF;
			14'd15091: ff_rdata <= 8'hFF;
			14'd15092: ff_rdata <= 8'hFF;
			14'd15093: ff_rdata <= 8'hFF;
			14'd15094: ff_rdata <= 8'hFF;
			14'd15095: ff_rdata <= 8'hFF;
			14'd15096: ff_rdata <= 8'hFF;
			14'd15097: ff_rdata <= 8'hFF;
			14'd15098: ff_rdata <= 8'hFF;
			14'd15099: ff_rdata <= 8'hFF;
			14'd15100: ff_rdata <= 8'hFF;
			14'd15101: ff_rdata <= 8'hFF;
			14'd15102: ff_rdata <= 8'hFF;
			14'd15103: ff_rdata <= 8'hFF;
			14'd15104: ff_rdata <= 8'hFF;
			14'd15105: ff_rdata <= 8'hFF;
			14'd15106: ff_rdata <= 8'hFF;
			14'd15107: ff_rdata <= 8'hFF;
			14'd15108: ff_rdata <= 8'hFF;
			14'd15109: ff_rdata <= 8'hFF;
			14'd15110: ff_rdata <= 8'hFF;
			14'd15111: ff_rdata <= 8'hFF;
			14'd15112: ff_rdata <= 8'hFF;
			14'd15113: ff_rdata <= 8'hFF;
			14'd15114: ff_rdata <= 8'hFF;
			14'd15115: ff_rdata <= 8'hFF;
			14'd15116: ff_rdata <= 8'hFF;
			14'd15117: ff_rdata <= 8'hFF;
			14'd15118: ff_rdata <= 8'hFF;
			14'd15119: ff_rdata <= 8'hFF;
			14'd15120: ff_rdata <= 8'hFF;
			14'd15121: ff_rdata <= 8'hFF;
			14'd15122: ff_rdata <= 8'hFF;
			14'd15123: ff_rdata <= 8'hFF;
			14'd15124: ff_rdata <= 8'hFF;
			14'd15125: ff_rdata <= 8'hFF;
			14'd15126: ff_rdata <= 8'hFF;
			14'd15127: ff_rdata <= 8'hFF;
			14'd15128: ff_rdata <= 8'hFF;
			14'd15129: ff_rdata <= 8'hFF;
			14'd15130: ff_rdata <= 8'hFF;
			14'd15131: ff_rdata <= 8'hFF;
			14'd15132: ff_rdata <= 8'hFF;
			14'd15133: ff_rdata <= 8'hFF;
			14'd15134: ff_rdata <= 8'hFF;
			14'd15135: ff_rdata <= 8'hFF;
			14'd15136: ff_rdata <= 8'hFF;
			14'd15137: ff_rdata <= 8'hFF;
			14'd15138: ff_rdata <= 8'hFF;
			14'd15139: ff_rdata <= 8'hFF;
			14'd15140: ff_rdata <= 8'hFF;
			14'd15141: ff_rdata <= 8'hFF;
			14'd15142: ff_rdata <= 8'hFF;
			14'd15143: ff_rdata <= 8'hFF;
			14'd15144: ff_rdata <= 8'hFF;
			14'd15145: ff_rdata <= 8'hFF;
			14'd15146: ff_rdata <= 8'hFF;
			14'd15147: ff_rdata <= 8'hFF;
			14'd15148: ff_rdata <= 8'hFF;
			14'd15149: ff_rdata <= 8'hFF;
			14'd15150: ff_rdata <= 8'hFF;
			14'd15151: ff_rdata <= 8'hFF;
			14'd15152: ff_rdata <= 8'hFF;
			14'd15153: ff_rdata <= 8'hFF;
			14'd15154: ff_rdata <= 8'hFF;
			14'd15155: ff_rdata <= 8'hFF;
			14'd15156: ff_rdata <= 8'hFF;
			14'd15157: ff_rdata <= 8'hFF;
			14'd15158: ff_rdata <= 8'hFF;
			14'd15159: ff_rdata <= 8'hFF;
			14'd15160: ff_rdata <= 8'hFF;
			14'd15161: ff_rdata <= 8'hFF;
			14'd15162: ff_rdata <= 8'hFF;
			14'd15163: ff_rdata <= 8'hFF;
			14'd15164: ff_rdata <= 8'hFF;
			14'd15165: ff_rdata <= 8'hFF;
			14'd15166: ff_rdata <= 8'hFF;
			14'd15167: ff_rdata <= 8'hFF;
			14'd15168: ff_rdata <= 8'hFF;
			14'd15169: ff_rdata <= 8'hFF;
			14'd15170: ff_rdata <= 8'hFF;
			14'd15171: ff_rdata <= 8'hFF;
			14'd15172: ff_rdata <= 8'hFF;
			14'd15173: ff_rdata <= 8'hFF;
			14'd15174: ff_rdata <= 8'hFF;
			14'd15175: ff_rdata <= 8'hFF;
			14'd15176: ff_rdata <= 8'hFF;
			14'd15177: ff_rdata <= 8'hFF;
			14'd15178: ff_rdata <= 8'hFF;
			14'd15179: ff_rdata <= 8'hFF;
			14'd15180: ff_rdata <= 8'hFF;
			14'd15181: ff_rdata <= 8'hFF;
			14'd15182: ff_rdata <= 8'hFF;
			14'd15183: ff_rdata <= 8'hFF;
			14'd15184: ff_rdata <= 8'hFF;
			14'd15185: ff_rdata <= 8'hFF;
			14'd15186: ff_rdata <= 8'hFF;
			14'd15187: ff_rdata <= 8'hFF;
			14'd15188: ff_rdata <= 8'hFF;
			14'd15189: ff_rdata <= 8'hFF;
			14'd15190: ff_rdata <= 8'hFF;
			14'd15191: ff_rdata <= 8'hFF;
			14'd15192: ff_rdata <= 8'hFF;
			14'd15193: ff_rdata <= 8'hFF;
			14'd15194: ff_rdata <= 8'hFF;
			14'd15195: ff_rdata <= 8'hFF;
			14'd15196: ff_rdata <= 8'hFF;
			14'd15197: ff_rdata <= 8'hFF;
			14'd15198: ff_rdata <= 8'hFF;
			14'd15199: ff_rdata <= 8'hFF;
			14'd15200: ff_rdata <= 8'hFF;
			14'd15201: ff_rdata <= 8'hFF;
			14'd15202: ff_rdata <= 8'hFF;
			14'd15203: ff_rdata <= 8'hFF;
			14'd15204: ff_rdata <= 8'hFF;
			14'd15205: ff_rdata <= 8'hFF;
			14'd15206: ff_rdata <= 8'hFF;
			14'd15207: ff_rdata <= 8'hFF;
			14'd15208: ff_rdata <= 8'hFF;
			14'd15209: ff_rdata <= 8'hFF;
			14'd15210: ff_rdata <= 8'hFF;
			14'd15211: ff_rdata <= 8'hFF;
			14'd15212: ff_rdata <= 8'hFF;
			14'd15213: ff_rdata <= 8'hFF;
			14'd15214: ff_rdata <= 8'hFF;
			14'd15215: ff_rdata <= 8'hFF;
			14'd15216: ff_rdata <= 8'hFF;
			14'd15217: ff_rdata <= 8'hFF;
			14'd15218: ff_rdata <= 8'hFF;
			14'd15219: ff_rdata <= 8'hFF;
			14'd15220: ff_rdata <= 8'hFF;
			14'd15221: ff_rdata <= 8'hFF;
			14'd15222: ff_rdata <= 8'hFF;
			14'd15223: ff_rdata <= 8'hFF;
			14'd15224: ff_rdata <= 8'hFF;
			14'd15225: ff_rdata <= 8'hFF;
			14'd15226: ff_rdata <= 8'hFF;
			14'd15227: ff_rdata <= 8'hFF;
			14'd15228: ff_rdata <= 8'hFF;
			14'd15229: ff_rdata <= 8'hFF;
			14'd15230: ff_rdata <= 8'hFF;
			14'd15231: ff_rdata <= 8'hFF;
			14'd15232: ff_rdata <= 8'hFF;
			14'd15233: ff_rdata <= 8'hFF;
			14'd15234: ff_rdata <= 8'hFF;
			14'd15235: ff_rdata <= 8'hFF;
			14'd15236: ff_rdata <= 8'hFF;
			14'd15237: ff_rdata <= 8'hFF;
			14'd15238: ff_rdata <= 8'hFF;
			14'd15239: ff_rdata <= 8'hFF;
			14'd15240: ff_rdata <= 8'hFF;
			14'd15241: ff_rdata <= 8'hFF;
			14'd15242: ff_rdata <= 8'hFF;
			14'd15243: ff_rdata <= 8'hFF;
			14'd15244: ff_rdata <= 8'hFF;
			14'd15245: ff_rdata <= 8'hFF;
			14'd15246: ff_rdata <= 8'hFF;
			14'd15247: ff_rdata <= 8'hFF;
			14'd15248: ff_rdata <= 8'hFF;
			14'd15249: ff_rdata <= 8'hFF;
			14'd15250: ff_rdata <= 8'hFF;
			14'd15251: ff_rdata <= 8'hFF;
			14'd15252: ff_rdata <= 8'hFF;
			14'd15253: ff_rdata <= 8'hFF;
			14'd15254: ff_rdata <= 8'hFF;
			14'd15255: ff_rdata <= 8'hFF;
			14'd15256: ff_rdata <= 8'hFF;
			14'd15257: ff_rdata <= 8'hFF;
			14'd15258: ff_rdata <= 8'hFF;
			14'd15259: ff_rdata <= 8'hFF;
			14'd15260: ff_rdata <= 8'hFF;
			14'd15261: ff_rdata <= 8'hFF;
			14'd15262: ff_rdata <= 8'hFF;
			14'd15263: ff_rdata <= 8'hFF;
			14'd15264: ff_rdata <= 8'hFF;
			14'd15265: ff_rdata <= 8'hFF;
			14'd15266: ff_rdata <= 8'hFF;
			14'd15267: ff_rdata <= 8'hFF;
			14'd15268: ff_rdata <= 8'hFF;
			14'd15269: ff_rdata <= 8'hFF;
			14'd15270: ff_rdata <= 8'hFF;
			14'd15271: ff_rdata <= 8'hFF;
			14'd15272: ff_rdata <= 8'hFF;
			14'd15273: ff_rdata <= 8'hFF;
			14'd15274: ff_rdata <= 8'hFF;
			14'd15275: ff_rdata <= 8'hFF;
			14'd15276: ff_rdata <= 8'hFF;
			14'd15277: ff_rdata <= 8'hFF;
			14'd15278: ff_rdata <= 8'hFF;
			14'd15279: ff_rdata <= 8'hFF;
			14'd15280: ff_rdata <= 8'hFF;
			14'd15281: ff_rdata <= 8'hFF;
			14'd15282: ff_rdata <= 8'hFF;
			14'd15283: ff_rdata <= 8'hFF;
			14'd15284: ff_rdata <= 8'hFF;
			14'd15285: ff_rdata <= 8'hFF;
			14'd15286: ff_rdata <= 8'hFF;
			14'd15287: ff_rdata <= 8'hFF;
			14'd15288: ff_rdata <= 8'hFF;
			14'd15289: ff_rdata <= 8'hFF;
			14'd15290: ff_rdata <= 8'hFF;
			14'd15291: ff_rdata <= 8'hFF;
			14'd15292: ff_rdata <= 8'hFF;
			14'd15293: ff_rdata <= 8'hFF;
			14'd15294: ff_rdata <= 8'hFF;
			14'd15295: ff_rdata <= 8'hFF;
			14'd15296: ff_rdata <= 8'hFF;
			14'd15297: ff_rdata <= 8'hFF;
			14'd15298: ff_rdata <= 8'hFF;
			14'd15299: ff_rdata <= 8'hFF;
			14'd15300: ff_rdata <= 8'hFF;
			14'd15301: ff_rdata <= 8'hFF;
			14'd15302: ff_rdata <= 8'hFF;
			14'd15303: ff_rdata <= 8'hFF;
			14'd15304: ff_rdata <= 8'hFF;
			14'd15305: ff_rdata <= 8'hFF;
			14'd15306: ff_rdata <= 8'hFF;
			14'd15307: ff_rdata <= 8'hFF;
			14'd15308: ff_rdata <= 8'hFF;
			14'd15309: ff_rdata <= 8'hFF;
			14'd15310: ff_rdata <= 8'hFF;
			14'd15311: ff_rdata <= 8'hFF;
			14'd15312: ff_rdata <= 8'hFF;
			14'd15313: ff_rdata <= 8'hFF;
			14'd15314: ff_rdata <= 8'hFF;
			14'd15315: ff_rdata <= 8'hFF;
			14'd15316: ff_rdata <= 8'hFF;
			14'd15317: ff_rdata <= 8'hFF;
			14'd15318: ff_rdata <= 8'hFF;
			14'd15319: ff_rdata <= 8'hFF;
			14'd15320: ff_rdata <= 8'hFF;
			14'd15321: ff_rdata <= 8'hFF;
			14'd15322: ff_rdata <= 8'hFF;
			14'd15323: ff_rdata <= 8'hFF;
			14'd15324: ff_rdata <= 8'hFF;
			14'd15325: ff_rdata <= 8'hFF;
			14'd15326: ff_rdata <= 8'hFF;
			14'd15327: ff_rdata <= 8'hFF;
			14'd15328: ff_rdata <= 8'hFF;
			14'd15329: ff_rdata <= 8'hFF;
			14'd15330: ff_rdata <= 8'hFF;
			14'd15331: ff_rdata <= 8'hFF;
			14'd15332: ff_rdata <= 8'hFF;
			14'd15333: ff_rdata <= 8'hFF;
			14'd15334: ff_rdata <= 8'hFF;
			14'd15335: ff_rdata <= 8'hFF;
			14'd15336: ff_rdata <= 8'hFF;
			14'd15337: ff_rdata <= 8'hFF;
			14'd15338: ff_rdata <= 8'hFF;
			14'd15339: ff_rdata <= 8'hFF;
			14'd15340: ff_rdata <= 8'hFF;
			14'd15341: ff_rdata <= 8'hFF;
			14'd15342: ff_rdata <= 8'hFF;
			14'd15343: ff_rdata <= 8'hFF;
			14'd15344: ff_rdata <= 8'hFF;
			14'd15345: ff_rdata <= 8'hFF;
			14'd15346: ff_rdata <= 8'hFF;
			14'd15347: ff_rdata <= 8'hFF;
			14'd15348: ff_rdata <= 8'hFF;
			14'd15349: ff_rdata <= 8'hFF;
			14'd15350: ff_rdata <= 8'hFF;
			14'd15351: ff_rdata <= 8'hFF;
			14'd15352: ff_rdata <= 8'hFF;
			14'd15353: ff_rdata <= 8'hFF;
			14'd15354: ff_rdata <= 8'hFF;
			14'd15355: ff_rdata <= 8'hFF;
			14'd15356: ff_rdata <= 8'hFF;
			14'd15357: ff_rdata <= 8'hFF;
			14'd15358: ff_rdata <= 8'hFF;
			14'd15359: ff_rdata <= 8'hFF;
			14'd15360: ff_rdata <= 8'hFF;
			14'd15361: ff_rdata <= 8'hFF;
			14'd15362: ff_rdata <= 8'hFF;
			14'd15363: ff_rdata <= 8'hFF;
			14'd15364: ff_rdata <= 8'hFF;
			14'd15365: ff_rdata <= 8'hFF;
			14'd15366: ff_rdata <= 8'hFF;
			14'd15367: ff_rdata <= 8'hFF;
			14'd15368: ff_rdata <= 8'hFF;
			14'd15369: ff_rdata <= 8'hFF;
			14'd15370: ff_rdata <= 8'hFF;
			14'd15371: ff_rdata <= 8'hFF;
			14'd15372: ff_rdata <= 8'hFF;
			14'd15373: ff_rdata <= 8'hFF;
			14'd15374: ff_rdata <= 8'hFF;
			14'd15375: ff_rdata <= 8'hFF;
			14'd15376: ff_rdata <= 8'hFF;
			14'd15377: ff_rdata <= 8'hFF;
			14'd15378: ff_rdata <= 8'hFF;
			14'd15379: ff_rdata <= 8'hFF;
			14'd15380: ff_rdata <= 8'hFF;
			14'd15381: ff_rdata <= 8'hFF;
			14'd15382: ff_rdata <= 8'hFF;
			14'd15383: ff_rdata <= 8'hFF;
			14'd15384: ff_rdata <= 8'hFF;
			14'd15385: ff_rdata <= 8'hFF;
			14'd15386: ff_rdata <= 8'hFF;
			14'd15387: ff_rdata <= 8'hFF;
			14'd15388: ff_rdata <= 8'hFF;
			14'd15389: ff_rdata <= 8'hFF;
			14'd15390: ff_rdata <= 8'hFF;
			14'd15391: ff_rdata <= 8'hFF;
			14'd15392: ff_rdata <= 8'hFF;
			14'd15393: ff_rdata <= 8'hFF;
			14'd15394: ff_rdata <= 8'hFF;
			14'd15395: ff_rdata <= 8'hFF;
			14'd15396: ff_rdata <= 8'hFF;
			14'd15397: ff_rdata <= 8'hFF;
			14'd15398: ff_rdata <= 8'hFF;
			14'd15399: ff_rdata <= 8'hFF;
			14'd15400: ff_rdata <= 8'hFF;
			14'd15401: ff_rdata <= 8'hFF;
			14'd15402: ff_rdata <= 8'hFF;
			14'd15403: ff_rdata <= 8'hFF;
			14'd15404: ff_rdata <= 8'hFF;
			14'd15405: ff_rdata <= 8'hFF;
			14'd15406: ff_rdata <= 8'hFF;
			14'd15407: ff_rdata <= 8'hFF;
			14'd15408: ff_rdata <= 8'hFF;
			14'd15409: ff_rdata <= 8'hFF;
			14'd15410: ff_rdata <= 8'hFF;
			14'd15411: ff_rdata <= 8'hFF;
			14'd15412: ff_rdata <= 8'hFF;
			14'd15413: ff_rdata <= 8'hFF;
			14'd15414: ff_rdata <= 8'hFF;
			14'd15415: ff_rdata <= 8'hFF;
			14'd15416: ff_rdata <= 8'hFF;
			14'd15417: ff_rdata <= 8'hFF;
			14'd15418: ff_rdata <= 8'hFF;
			14'd15419: ff_rdata <= 8'hFF;
			14'd15420: ff_rdata <= 8'hFF;
			14'd15421: ff_rdata <= 8'hFF;
			14'd15422: ff_rdata <= 8'hFF;
			14'd15423: ff_rdata <= 8'hFF;
			14'd15424: ff_rdata <= 8'hFF;
			14'd15425: ff_rdata <= 8'hFF;
			14'd15426: ff_rdata <= 8'hFF;
			14'd15427: ff_rdata <= 8'hFF;
			14'd15428: ff_rdata <= 8'hFF;
			14'd15429: ff_rdata <= 8'hFF;
			14'd15430: ff_rdata <= 8'hFF;
			14'd15431: ff_rdata <= 8'hFF;
			14'd15432: ff_rdata <= 8'hFF;
			14'd15433: ff_rdata <= 8'hFF;
			14'd15434: ff_rdata <= 8'hFF;
			14'd15435: ff_rdata <= 8'hFF;
			14'd15436: ff_rdata <= 8'hFF;
			14'd15437: ff_rdata <= 8'hFF;
			14'd15438: ff_rdata <= 8'hFF;
			14'd15439: ff_rdata <= 8'hFF;
			14'd15440: ff_rdata <= 8'hFF;
			14'd15441: ff_rdata <= 8'hFF;
			14'd15442: ff_rdata <= 8'hFF;
			14'd15443: ff_rdata <= 8'hFF;
			14'd15444: ff_rdata <= 8'hFF;
			14'd15445: ff_rdata <= 8'hFF;
			14'd15446: ff_rdata <= 8'hFF;
			14'd15447: ff_rdata <= 8'hFF;
			14'd15448: ff_rdata <= 8'hFF;
			14'd15449: ff_rdata <= 8'hFF;
			14'd15450: ff_rdata <= 8'hFF;
			14'd15451: ff_rdata <= 8'hFF;
			14'd15452: ff_rdata <= 8'hFF;
			14'd15453: ff_rdata <= 8'hFF;
			14'd15454: ff_rdata <= 8'hFF;
			14'd15455: ff_rdata <= 8'hFF;
			14'd15456: ff_rdata <= 8'hFF;
			14'd15457: ff_rdata <= 8'hFF;
			14'd15458: ff_rdata <= 8'hFF;
			14'd15459: ff_rdata <= 8'hFF;
			14'd15460: ff_rdata <= 8'hFF;
			14'd15461: ff_rdata <= 8'hFF;
			14'd15462: ff_rdata <= 8'hFF;
			14'd15463: ff_rdata <= 8'hFF;
			14'd15464: ff_rdata <= 8'hFF;
			14'd15465: ff_rdata <= 8'hFF;
			14'd15466: ff_rdata <= 8'hFF;
			14'd15467: ff_rdata <= 8'hFF;
			14'd15468: ff_rdata <= 8'hFF;
			14'd15469: ff_rdata <= 8'hFF;
			14'd15470: ff_rdata <= 8'hFF;
			14'd15471: ff_rdata <= 8'hFF;
			14'd15472: ff_rdata <= 8'hFF;
			14'd15473: ff_rdata <= 8'hFF;
			14'd15474: ff_rdata <= 8'hFF;
			14'd15475: ff_rdata <= 8'hFF;
			14'd15476: ff_rdata <= 8'hFF;
			14'd15477: ff_rdata <= 8'hFF;
			14'd15478: ff_rdata <= 8'hFF;
			14'd15479: ff_rdata <= 8'hFF;
			14'd15480: ff_rdata <= 8'hFF;
			14'd15481: ff_rdata <= 8'hFF;
			14'd15482: ff_rdata <= 8'hFF;
			14'd15483: ff_rdata <= 8'hFF;
			14'd15484: ff_rdata <= 8'hFF;
			14'd15485: ff_rdata <= 8'hFF;
			14'd15486: ff_rdata <= 8'hFF;
			14'd15487: ff_rdata <= 8'hFF;
			14'd15488: ff_rdata <= 8'hFF;
			14'd15489: ff_rdata <= 8'hFF;
			14'd15490: ff_rdata <= 8'hFF;
			14'd15491: ff_rdata <= 8'hFF;
			14'd15492: ff_rdata <= 8'hFF;
			14'd15493: ff_rdata <= 8'hFF;
			14'd15494: ff_rdata <= 8'hFF;
			14'd15495: ff_rdata <= 8'hFF;
			14'd15496: ff_rdata <= 8'hFF;
			14'd15497: ff_rdata <= 8'hFF;
			14'd15498: ff_rdata <= 8'hFF;
			14'd15499: ff_rdata <= 8'hFF;
			14'd15500: ff_rdata <= 8'hFF;
			14'd15501: ff_rdata <= 8'hFF;
			14'd15502: ff_rdata <= 8'hFF;
			14'd15503: ff_rdata <= 8'hFF;
			14'd15504: ff_rdata <= 8'hFF;
			14'd15505: ff_rdata <= 8'hFF;
			14'd15506: ff_rdata <= 8'hFF;
			14'd15507: ff_rdata <= 8'hFF;
			14'd15508: ff_rdata <= 8'hFF;
			14'd15509: ff_rdata <= 8'hFF;
			14'd15510: ff_rdata <= 8'hFF;
			14'd15511: ff_rdata <= 8'hFF;
			14'd15512: ff_rdata <= 8'hFF;
			14'd15513: ff_rdata <= 8'hFF;
			14'd15514: ff_rdata <= 8'hFF;
			14'd15515: ff_rdata <= 8'hFF;
			14'd15516: ff_rdata <= 8'hFF;
			14'd15517: ff_rdata <= 8'hFF;
			14'd15518: ff_rdata <= 8'hFF;
			14'd15519: ff_rdata <= 8'hFF;
			14'd15520: ff_rdata <= 8'hFF;
			14'd15521: ff_rdata <= 8'hFF;
			14'd15522: ff_rdata <= 8'hFF;
			14'd15523: ff_rdata <= 8'hFF;
			14'd15524: ff_rdata <= 8'hFF;
			14'd15525: ff_rdata <= 8'hFF;
			14'd15526: ff_rdata <= 8'hFF;
			14'd15527: ff_rdata <= 8'hFF;
			14'd15528: ff_rdata <= 8'hFF;
			14'd15529: ff_rdata <= 8'hFF;
			14'd15530: ff_rdata <= 8'hFF;
			14'd15531: ff_rdata <= 8'hFF;
			14'd15532: ff_rdata <= 8'hFF;
			14'd15533: ff_rdata <= 8'hFF;
			14'd15534: ff_rdata <= 8'hFF;
			14'd15535: ff_rdata <= 8'hFF;
			14'd15536: ff_rdata <= 8'hFF;
			14'd15537: ff_rdata <= 8'hFF;
			14'd15538: ff_rdata <= 8'hFF;
			14'd15539: ff_rdata <= 8'hFF;
			14'd15540: ff_rdata <= 8'hFF;
			14'd15541: ff_rdata <= 8'hFF;
			14'd15542: ff_rdata <= 8'hFF;
			14'd15543: ff_rdata <= 8'hFF;
			14'd15544: ff_rdata <= 8'hFF;
			14'd15545: ff_rdata <= 8'hFF;
			14'd15546: ff_rdata <= 8'hFF;
			14'd15547: ff_rdata <= 8'hFF;
			14'd15548: ff_rdata <= 8'hFF;
			14'd15549: ff_rdata <= 8'hFF;
			14'd15550: ff_rdata <= 8'hFF;
			14'd15551: ff_rdata <= 8'hFF;
			14'd15552: ff_rdata <= 8'hFF;
			14'd15553: ff_rdata <= 8'hFF;
			14'd15554: ff_rdata <= 8'hFF;
			14'd15555: ff_rdata <= 8'hFF;
			14'd15556: ff_rdata <= 8'hFF;
			14'd15557: ff_rdata <= 8'hFF;
			14'd15558: ff_rdata <= 8'hFF;
			14'd15559: ff_rdata <= 8'hFF;
			14'd15560: ff_rdata <= 8'hFF;
			14'd15561: ff_rdata <= 8'hFF;
			14'd15562: ff_rdata <= 8'hFF;
			14'd15563: ff_rdata <= 8'hFF;
			14'd15564: ff_rdata <= 8'hFF;
			14'd15565: ff_rdata <= 8'hFF;
			14'd15566: ff_rdata <= 8'hFF;
			14'd15567: ff_rdata <= 8'hFF;
			14'd15568: ff_rdata <= 8'hFF;
			14'd15569: ff_rdata <= 8'hFF;
			14'd15570: ff_rdata <= 8'hFF;
			14'd15571: ff_rdata <= 8'hFF;
			14'd15572: ff_rdata <= 8'hFF;
			14'd15573: ff_rdata <= 8'hFF;
			14'd15574: ff_rdata <= 8'hFF;
			14'd15575: ff_rdata <= 8'hFF;
			14'd15576: ff_rdata <= 8'hFF;
			14'd15577: ff_rdata <= 8'hFF;
			14'd15578: ff_rdata <= 8'hFF;
			14'd15579: ff_rdata <= 8'hFF;
			14'd15580: ff_rdata <= 8'hFF;
			14'd15581: ff_rdata <= 8'hFF;
			14'd15582: ff_rdata <= 8'hFF;
			14'd15583: ff_rdata <= 8'hFF;
			14'd15584: ff_rdata <= 8'hFF;
			14'd15585: ff_rdata <= 8'hFF;
			14'd15586: ff_rdata <= 8'hFF;
			14'd15587: ff_rdata <= 8'hFF;
			14'd15588: ff_rdata <= 8'hFF;
			14'd15589: ff_rdata <= 8'hFF;
			14'd15590: ff_rdata <= 8'hFF;
			14'd15591: ff_rdata <= 8'hFF;
			14'd15592: ff_rdata <= 8'hFF;
			14'd15593: ff_rdata <= 8'hFF;
			14'd15594: ff_rdata <= 8'hFF;
			14'd15595: ff_rdata <= 8'hFF;
			14'd15596: ff_rdata <= 8'hFF;
			14'd15597: ff_rdata <= 8'hFF;
			14'd15598: ff_rdata <= 8'hFF;
			14'd15599: ff_rdata <= 8'hFF;
			14'd15600: ff_rdata <= 8'hFF;
			14'd15601: ff_rdata <= 8'hFF;
			14'd15602: ff_rdata <= 8'hFF;
			14'd15603: ff_rdata <= 8'hFF;
			14'd15604: ff_rdata <= 8'hFF;
			14'd15605: ff_rdata <= 8'hFF;
			14'd15606: ff_rdata <= 8'hFF;
			14'd15607: ff_rdata <= 8'hFF;
			14'd15608: ff_rdata <= 8'hFF;
			14'd15609: ff_rdata <= 8'hFF;
			14'd15610: ff_rdata <= 8'hFF;
			14'd15611: ff_rdata <= 8'hFF;
			14'd15612: ff_rdata <= 8'hFF;
			14'd15613: ff_rdata <= 8'hFF;
			14'd15614: ff_rdata <= 8'hFF;
			14'd15615: ff_rdata <= 8'hFF;
			14'd15616: ff_rdata <= 8'hFF;
			14'd15617: ff_rdata <= 8'hFF;
			14'd15618: ff_rdata <= 8'hFF;
			14'd15619: ff_rdata <= 8'hFF;
			14'd15620: ff_rdata <= 8'hFF;
			14'd15621: ff_rdata <= 8'hFF;
			14'd15622: ff_rdata <= 8'hFF;
			14'd15623: ff_rdata <= 8'hFF;
			14'd15624: ff_rdata <= 8'hFF;
			14'd15625: ff_rdata <= 8'hFF;
			14'd15626: ff_rdata <= 8'hFF;
			14'd15627: ff_rdata <= 8'hFF;
			14'd15628: ff_rdata <= 8'hFF;
			14'd15629: ff_rdata <= 8'hFF;
			14'd15630: ff_rdata <= 8'hFF;
			14'd15631: ff_rdata <= 8'hFF;
			14'd15632: ff_rdata <= 8'hFF;
			14'd15633: ff_rdata <= 8'hFF;
			14'd15634: ff_rdata <= 8'hFF;
			14'd15635: ff_rdata <= 8'hFF;
			14'd15636: ff_rdata <= 8'hFF;
			14'd15637: ff_rdata <= 8'hFF;
			14'd15638: ff_rdata <= 8'hFF;
			14'd15639: ff_rdata <= 8'hFF;
			14'd15640: ff_rdata <= 8'hFF;
			14'd15641: ff_rdata <= 8'hFF;
			14'd15642: ff_rdata <= 8'hFF;
			14'd15643: ff_rdata <= 8'hFF;
			14'd15644: ff_rdata <= 8'hFF;
			14'd15645: ff_rdata <= 8'hFF;
			14'd15646: ff_rdata <= 8'hFF;
			14'd15647: ff_rdata <= 8'hFF;
			14'd15648: ff_rdata <= 8'hFF;
			14'd15649: ff_rdata <= 8'hFF;
			14'd15650: ff_rdata <= 8'hFF;
			14'd15651: ff_rdata <= 8'hFF;
			14'd15652: ff_rdata <= 8'hFF;
			14'd15653: ff_rdata <= 8'hFF;
			14'd15654: ff_rdata <= 8'hFF;
			14'd15655: ff_rdata <= 8'hFF;
			14'd15656: ff_rdata <= 8'hFF;
			14'd15657: ff_rdata <= 8'hFF;
			14'd15658: ff_rdata <= 8'hFF;
			14'd15659: ff_rdata <= 8'hFF;
			14'd15660: ff_rdata <= 8'hFF;
			14'd15661: ff_rdata <= 8'hFF;
			14'd15662: ff_rdata <= 8'hFF;
			14'd15663: ff_rdata <= 8'hFF;
			14'd15664: ff_rdata <= 8'hFF;
			14'd15665: ff_rdata <= 8'hFF;
			14'd15666: ff_rdata <= 8'hFF;
			14'd15667: ff_rdata <= 8'hFF;
			14'd15668: ff_rdata <= 8'hFF;
			14'd15669: ff_rdata <= 8'hFF;
			14'd15670: ff_rdata <= 8'hFF;
			14'd15671: ff_rdata <= 8'hFF;
			14'd15672: ff_rdata <= 8'hFF;
			14'd15673: ff_rdata <= 8'hFF;
			14'd15674: ff_rdata <= 8'hFF;
			14'd15675: ff_rdata <= 8'hFF;
			14'd15676: ff_rdata <= 8'hFF;
			14'd15677: ff_rdata <= 8'hFF;
			14'd15678: ff_rdata <= 8'hFF;
			14'd15679: ff_rdata <= 8'hFF;
			14'd15680: ff_rdata <= 8'hFF;
			14'd15681: ff_rdata <= 8'hFF;
			14'd15682: ff_rdata <= 8'hFF;
			14'd15683: ff_rdata <= 8'hFF;
			14'd15684: ff_rdata <= 8'hFF;
			14'd15685: ff_rdata <= 8'hFF;
			14'd15686: ff_rdata <= 8'hFF;
			14'd15687: ff_rdata <= 8'hFF;
			14'd15688: ff_rdata <= 8'hFF;
			14'd15689: ff_rdata <= 8'hFF;
			14'd15690: ff_rdata <= 8'hFF;
			14'd15691: ff_rdata <= 8'hFF;
			14'd15692: ff_rdata <= 8'hFF;
			14'd15693: ff_rdata <= 8'hFF;
			14'd15694: ff_rdata <= 8'hFF;
			14'd15695: ff_rdata <= 8'hFF;
			14'd15696: ff_rdata <= 8'hFF;
			14'd15697: ff_rdata <= 8'hFF;
			14'd15698: ff_rdata <= 8'hFF;
			14'd15699: ff_rdata <= 8'hFF;
			14'd15700: ff_rdata <= 8'hFF;
			14'd15701: ff_rdata <= 8'hFF;
			14'd15702: ff_rdata <= 8'hFF;
			14'd15703: ff_rdata <= 8'hFF;
			14'd15704: ff_rdata <= 8'hFF;
			14'd15705: ff_rdata <= 8'hFF;
			14'd15706: ff_rdata <= 8'hFF;
			14'd15707: ff_rdata <= 8'hFF;
			14'd15708: ff_rdata <= 8'hFF;
			14'd15709: ff_rdata <= 8'hFF;
			14'd15710: ff_rdata <= 8'hFF;
			14'd15711: ff_rdata <= 8'hFF;
			14'd15712: ff_rdata <= 8'hFF;
			14'd15713: ff_rdata <= 8'hFF;
			14'd15714: ff_rdata <= 8'hFF;
			14'd15715: ff_rdata <= 8'hFF;
			14'd15716: ff_rdata <= 8'hFF;
			14'd15717: ff_rdata <= 8'hFF;
			14'd15718: ff_rdata <= 8'hFF;
			14'd15719: ff_rdata <= 8'hFF;
			14'd15720: ff_rdata <= 8'hFF;
			14'd15721: ff_rdata <= 8'hFF;
			14'd15722: ff_rdata <= 8'hFF;
			14'd15723: ff_rdata <= 8'hFF;
			14'd15724: ff_rdata <= 8'hFF;
			14'd15725: ff_rdata <= 8'hFF;
			14'd15726: ff_rdata <= 8'hFF;
			14'd15727: ff_rdata <= 8'hFF;
			14'd15728: ff_rdata <= 8'hFF;
			14'd15729: ff_rdata <= 8'hFF;
			14'd15730: ff_rdata <= 8'hFF;
			14'd15731: ff_rdata <= 8'hFF;
			14'd15732: ff_rdata <= 8'hFF;
			14'd15733: ff_rdata <= 8'hFF;
			14'd15734: ff_rdata <= 8'hFF;
			14'd15735: ff_rdata <= 8'hFF;
			14'd15736: ff_rdata <= 8'hFF;
			14'd15737: ff_rdata <= 8'hFF;
			14'd15738: ff_rdata <= 8'hFF;
			14'd15739: ff_rdata <= 8'hFF;
			14'd15740: ff_rdata <= 8'hFF;
			14'd15741: ff_rdata <= 8'hFF;
			14'd15742: ff_rdata <= 8'hFF;
			14'd15743: ff_rdata <= 8'hFF;
			14'd15744: ff_rdata <= 8'hFF;
			14'd15745: ff_rdata <= 8'hFF;
			14'd15746: ff_rdata <= 8'hFF;
			14'd15747: ff_rdata <= 8'hFF;
			14'd15748: ff_rdata <= 8'hFF;
			14'd15749: ff_rdata <= 8'hFF;
			14'd15750: ff_rdata <= 8'hFF;
			14'd15751: ff_rdata <= 8'hFF;
			14'd15752: ff_rdata <= 8'hFF;
			14'd15753: ff_rdata <= 8'hFF;
			14'd15754: ff_rdata <= 8'hFF;
			14'd15755: ff_rdata <= 8'hFF;
			14'd15756: ff_rdata <= 8'hFF;
			14'd15757: ff_rdata <= 8'hFF;
			14'd15758: ff_rdata <= 8'hFF;
			14'd15759: ff_rdata <= 8'hFF;
			14'd15760: ff_rdata <= 8'hFF;
			14'd15761: ff_rdata <= 8'hFF;
			14'd15762: ff_rdata <= 8'hFF;
			14'd15763: ff_rdata <= 8'hFF;
			14'd15764: ff_rdata <= 8'hFF;
			14'd15765: ff_rdata <= 8'hFF;
			14'd15766: ff_rdata <= 8'hFF;
			14'd15767: ff_rdata <= 8'hFF;
			14'd15768: ff_rdata <= 8'hFF;
			14'd15769: ff_rdata <= 8'hFF;
			14'd15770: ff_rdata <= 8'hFF;
			14'd15771: ff_rdata <= 8'hFF;
			14'd15772: ff_rdata <= 8'hFF;
			14'd15773: ff_rdata <= 8'hFF;
			14'd15774: ff_rdata <= 8'hFF;
			14'd15775: ff_rdata <= 8'hFF;
			14'd15776: ff_rdata <= 8'hFF;
			14'd15777: ff_rdata <= 8'hFF;
			14'd15778: ff_rdata <= 8'hFF;
			14'd15779: ff_rdata <= 8'hFF;
			14'd15780: ff_rdata <= 8'hFF;
			14'd15781: ff_rdata <= 8'hFF;
			14'd15782: ff_rdata <= 8'hFF;
			14'd15783: ff_rdata <= 8'hFF;
			14'd15784: ff_rdata <= 8'hFF;
			14'd15785: ff_rdata <= 8'hFF;
			14'd15786: ff_rdata <= 8'hFF;
			14'd15787: ff_rdata <= 8'hFF;
			14'd15788: ff_rdata <= 8'hFF;
			14'd15789: ff_rdata <= 8'hFF;
			14'd15790: ff_rdata <= 8'hFF;
			14'd15791: ff_rdata <= 8'hFF;
			14'd15792: ff_rdata <= 8'hFF;
			14'd15793: ff_rdata <= 8'hFF;
			14'd15794: ff_rdata <= 8'hFF;
			14'd15795: ff_rdata <= 8'hFF;
			14'd15796: ff_rdata <= 8'hFF;
			14'd15797: ff_rdata <= 8'hFF;
			14'd15798: ff_rdata <= 8'hFF;
			14'd15799: ff_rdata <= 8'hFF;
			14'd15800: ff_rdata <= 8'hFF;
			14'd15801: ff_rdata <= 8'hFF;
			14'd15802: ff_rdata <= 8'hFF;
			14'd15803: ff_rdata <= 8'hFF;
			14'd15804: ff_rdata <= 8'hFF;
			14'd15805: ff_rdata <= 8'hFF;
			14'd15806: ff_rdata <= 8'hFF;
			14'd15807: ff_rdata <= 8'hFF;
			14'd15808: ff_rdata <= 8'hFF;
			14'd15809: ff_rdata <= 8'hFF;
			14'd15810: ff_rdata <= 8'hFF;
			14'd15811: ff_rdata <= 8'hFF;
			14'd15812: ff_rdata <= 8'hFF;
			14'd15813: ff_rdata <= 8'hFF;
			14'd15814: ff_rdata <= 8'hFF;
			14'd15815: ff_rdata <= 8'hFF;
			14'd15816: ff_rdata <= 8'hFF;
			14'd15817: ff_rdata <= 8'hFF;
			14'd15818: ff_rdata <= 8'hFF;
			14'd15819: ff_rdata <= 8'hFF;
			14'd15820: ff_rdata <= 8'hFF;
			14'd15821: ff_rdata <= 8'hFF;
			14'd15822: ff_rdata <= 8'hFF;
			14'd15823: ff_rdata <= 8'hFF;
			14'd15824: ff_rdata <= 8'hFF;
			14'd15825: ff_rdata <= 8'hFF;
			14'd15826: ff_rdata <= 8'hFF;
			14'd15827: ff_rdata <= 8'hFF;
			14'd15828: ff_rdata <= 8'hFF;
			14'd15829: ff_rdata <= 8'hFF;
			14'd15830: ff_rdata <= 8'hFF;
			14'd15831: ff_rdata <= 8'hFF;
			14'd15832: ff_rdata <= 8'hFF;
			14'd15833: ff_rdata <= 8'hFF;
			14'd15834: ff_rdata <= 8'hFF;
			14'd15835: ff_rdata <= 8'hFF;
			14'd15836: ff_rdata <= 8'hFF;
			14'd15837: ff_rdata <= 8'hFF;
			14'd15838: ff_rdata <= 8'hFF;
			14'd15839: ff_rdata <= 8'hFF;
			14'd15840: ff_rdata <= 8'hFF;
			14'd15841: ff_rdata <= 8'hFF;
			14'd15842: ff_rdata <= 8'hFF;
			14'd15843: ff_rdata <= 8'hFF;
			14'd15844: ff_rdata <= 8'hFF;
			14'd15845: ff_rdata <= 8'hFF;
			14'd15846: ff_rdata <= 8'hFF;
			14'd15847: ff_rdata <= 8'hFF;
			14'd15848: ff_rdata <= 8'hFF;
			14'd15849: ff_rdata <= 8'hFF;
			14'd15850: ff_rdata <= 8'hFF;
			14'd15851: ff_rdata <= 8'hFF;
			14'd15852: ff_rdata <= 8'hFF;
			14'd15853: ff_rdata <= 8'hFF;
			14'd15854: ff_rdata <= 8'hFF;
			14'd15855: ff_rdata <= 8'hFF;
			14'd15856: ff_rdata <= 8'hFF;
			14'd15857: ff_rdata <= 8'hFF;
			14'd15858: ff_rdata <= 8'hFF;
			14'd15859: ff_rdata <= 8'hFF;
			14'd15860: ff_rdata <= 8'hFF;
			14'd15861: ff_rdata <= 8'hFF;
			14'd15862: ff_rdata <= 8'hFF;
			14'd15863: ff_rdata <= 8'hFF;
			14'd15864: ff_rdata <= 8'hFF;
			14'd15865: ff_rdata <= 8'hFF;
			14'd15866: ff_rdata <= 8'hFF;
			14'd15867: ff_rdata <= 8'hFF;
			14'd15868: ff_rdata <= 8'hFF;
			14'd15869: ff_rdata <= 8'hFF;
			14'd15870: ff_rdata <= 8'hFF;
			14'd15871: ff_rdata <= 8'hFF;
			14'd15872: ff_rdata <= 8'hFF;
			14'd15873: ff_rdata <= 8'hFF;
			14'd15874: ff_rdata <= 8'hFF;
			14'd15875: ff_rdata <= 8'hFF;
			14'd15876: ff_rdata <= 8'hFF;
			14'd15877: ff_rdata <= 8'hFF;
			14'd15878: ff_rdata <= 8'hFF;
			14'd15879: ff_rdata <= 8'hFF;
			14'd15880: ff_rdata <= 8'hFF;
			14'd15881: ff_rdata <= 8'hFF;
			14'd15882: ff_rdata <= 8'hFF;
			14'd15883: ff_rdata <= 8'hFF;
			14'd15884: ff_rdata <= 8'hFF;
			14'd15885: ff_rdata <= 8'hFF;
			14'd15886: ff_rdata <= 8'hFF;
			14'd15887: ff_rdata <= 8'hFF;
			14'd15888: ff_rdata <= 8'hFF;
			14'd15889: ff_rdata <= 8'hFF;
			14'd15890: ff_rdata <= 8'hFF;
			14'd15891: ff_rdata <= 8'hFF;
			14'd15892: ff_rdata <= 8'hFF;
			14'd15893: ff_rdata <= 8'hFF;
			14'd15894: ff_rdata <= 8'hFF;
			14'd15895: ff_rdata <= 8'hFF;
			14'd15896: ff_rdata <= 8'hFF;
			14'd15897: ff_rdata <= 8'hFF;
			14'd15898: ff_rdata <= 8'hFF;
			14'd15899: ff_rdata <= 8'hFF;
			14'd15900: ff_rdata <= 8'hFF;
			14'd15901: ff_rdata <= 8'hFF;
			14'd15902: ff_rdata <= 8'hFF;
			14'd15903: ff_rdata <= 8'hFF;
			14'd15904: ff_rdata <= 8'hFF;
			14'd15905: ff_rdata <= 8'hFF;
			14'd15906: ff_rdata <= 8'hFF;
			14'd15907: ff_rdata <= 8'hFF;
			14'd15908: ff_rdata <= 8'hFF;
			14'd15909: ff_rdata <= 8'hFF;
			14'd15910: ff_rdata <= 8'hFF;
			14'd15911: ff_rdata <= 8'hFF;
			14'd15912: ff_rdata <= 8'hFF;
			14'd15913: ff_rdata <= 8'hFF;
			14'd15914: ff_rdata <= 8'hFF;
			14'd15915: ff_rdata <= 8'hFF;
			14'd15916: ff_rdata <= 8'hFF;
			14'd15917: ff_rdata <= 8'hFF;
			14'd15918: ff_rdata <= 8'hFF;
			14'd15919: ff_rdata <= 8'hFF;
			14'd15920: ff_rdata <= 8'hFF;
			14'd15921: ff_rdata <= 8'hFF;
			14'd15922: ff_rdata <= 8'hFF;
			14'd15923: ff_rdata <= 8'hFF;
			14'd15924: ff_rdata <= 8'hFF;
			14'd15925: ff_rdata <= 8'hFF;
			14'd15926: ff_rdata <= 8'hFF;
			14'd15927: ff_rdata <= 8'hFF;
			14'd15928: ff_rdata <= 8'hFF;
			14'd15929: ff_rdata <= 8'hFF;
			14'd15930: ff_rdata <= 8'hFF;
			14'd15931: ff_rdata <= 8'hFF;
			14'd15932: ff_rdata <= 8'hFF;
			14'd15933: ff_rdata <= 8'hFF;
			14'd15934: ff_rdata <= 8'hFF;
			14'd15935: ff_rdata <= 8'hFF;
			14'd15936: ff_rdata <= 8'hFF;
			14'd15937: ff_rdata <= 8'hFF;
			14'd15938: ff_rdata <= 8'hFF;
			14'd15939: ff_rdata <= 8'hFF;
			14'd15940: ff_rdata <= 8'hFF;
			14'd15941: ff_rdata <= 8'hFF;
			14'd15942: ff_rdata <= 8'hFF;
			14'd15943: ff_rdata <= 8'hFF;
			14'd15944: ff_rdata <= 8'hFF;
			14'd15945: ff_rdata <= 8'hFF;
			14'd15946: ff_rdata <= 8'hFF;
			14'd15947: ff_rdata <= 8'hFF;
			14'd15948: ff_rdata <= 8'hFF;
			14'd15949: ff_rdata <= 8'hFF;
			14'd15950: ff_rdata <= 8'hFF;
			14'd15951: ff_rdata <= 8'hFF;
			14'd15952: ff_rdata <= 8'hFF;
			14'd15953: ff_rdata <= 8'hFF;
			14'd15954: ff_rdata <= 8'hFF;
			14'd15955: ff_rdata <= 8'hFF;
			14'd15956: ff_rdata <= 8'hFF;
			14'd15957: ff_rdata <= 8'hFF;
			14'd15958: ff_rdata <= 8'hFF;
			14'd15959: ff_rdata <= 8'hFF;
			14'd15960: ff_rdata <= 8'hFF;
			14'd15961: ff_rdata <= 8'hFF;
			14'd15962: ff_rdata <= 8'hFF;
			14'd15963: ff_rdata <= 8'hFF;
			14'd15964: ff_rdata <= 8'hFF;
			14'd15965: ff_rdata <= 8'hFF;
			14'd15966: ff_rdata <= 8'hFF;
			14'd15967: ff_rdata <= 8'hFF;
			14'd15968: ff_rdata <= 8'hFF;
			14'd15969: ff_rdata <= 8'hFF;
			14'd15970: ff_rdata <= 8'hFF;
			14'd15971: ff_rdata <= 8'hFF;
			14'd15972: ff_rdata <= 8'hFF;
			14'd15973: ff_rdata <= 8'hFF;
			14'd15974: ff_rdata <= 8'hFF;
			14'd15975: ff_rdata <= 8'hFF;
			14'd15976: ff_rdata <= 8'hFF;
			14'd15977: ff_rdata <= 8'hFF;
			14'd15978: ff_rdata <= 8'hFF;
			14'd15979: ff_rdata <= 8'hFF;
			14'd15980: ff_rdata <= 8'hFF;
			14'd15981: ff_rdata <= 8'hFF;
			14'd15982: ff_rdata <= 8'hFF;
			14'd15983: ff_rdata <= 8'hFF;
			14'd15984: ff_rdata <= 8'hFF;
			14'd15985: ff_rdata <= 8'hFF;
			14'd15986: ff_rdata <= 8'hFF;
			14'd15987: ff_rdata <= 8'hFF;
			14'd15988: ff_rdata <= 8'hFF;
			14'd15989: ff_rdata <= 8'hFF;
			14'd15990: ff_rdata <= 8'hFF;
			14'd15991: ff_rdata <= 8'hFF;
			14'd15992: ff_rdata <= 8'hFF;
			14'd15993: ff_rdata <= 8'hFF;
			14'd15994: ff_rdata <= 8'hFF;
			14'd15995: ff_rdata <= 8'hFF;
			14'd15996: ff_rdata <= 8'hFF;
			14'd15997: ff_rdata <= 8'hFF;
			14'd15998: ff_rdata <= 8'hFF;
			14'd15999: ff_rdata <= 8'hFF;
			14'd16000: ff_rdata <= 8'hFF;
			14'd16001: ff_rdata <= 8'hFF;
			14'd16002: ff_rdata <= 8'hFF;
			14'd16003: ff_rdata <= 8'hFF;
			14'd16004: ff_rdata <= 8'hFF;
			14'd16005: ff_rdata <= 8'hFF;
			14'd16006: ff_rdata <= 8'hFF;
			14'd16007: ff_rdata <= 8'hFF;
			14'd16008: ff_rdata <= 8'hFF;
			14'd16009: ff_rdata <= 8'hFF;
			14'd16010: ff_rdata <= 8'hFF;
			14'd16011: ff_rdata <= 8'hFF;
			14'd16012: ff_rdata <= 8'hFF;
			14'd16013: ff_rdata <= 8'hFF;
			14'd16014: ff_rdata <= 8'hFF;
			14'd16015: ff_rdata <= 8'hFF;
			14'd16016: ff_rdata <= 8'hFF;
			14'd16017: ff_rdata <= 8'hFF;
			14'd16018: ff_rdata <= 8'hFF;
			14'd16019: ff_rdata <= 8'hFF;
			14'd16020: ff_rdata <= 8'hFF;
			14'd16021: ff_rdata <= 8'hFF;
			14'd16022: ff_rdata <= 8'hFF;
			14'd16023: ff_rdata <= 8'hFF;
			14'd16024: ff_rdata <= 8'hFF;
			14'd16025: ff_rdata <= 8'hFF;
			14'd16026: ff_rdata <= 8'hFF;
			14'd16027: ff_rdata <= 8'hFF;
			14'd16028: ff_rdata <= 8'hFF;
			14'd16029: ff_rdata <= 8'hFF;
			14'd16030: ff_rdata <= 8'hFF;
			14'd16031: ff_rdata <= 8'hFF;
			14'd16032: ff_rdata <= 8'hFF;
			14'd16033: ff_rdata <= 8'hFF;
			14'd16034: ff_rdata <= 8'hFF;
			14'd16035: ff_rdata <= 8'hFF;
			14'd16036: ff_rdata <= 8'hFF;
			14'd16037: ff_rdata <= 8'hFF;
			14'd16038: ff_rdata <= 8'hFF;
			14'd16039: ff_rdata <= 8'hFF;
			14'd16040: ff_rdata <= 8'hFF;
			14'd16041: ff_rdata <= 8'hFF;
			14'd16042: ff_rdata <= 8'hFF;
			14'd16043: ff_rdata <= 8'hFF;
			14'd16044: ff_rdata <= 8'hFF;
			14'd16045: ff_rdata <= 8'hFF;
			14'd16046: ff_rdata <= 8'hFF;
			14'd16047: ff_rdata <= 8'hFF;
			14'd16048: ff_rdata <= 8'hFF;
			14'd16049: ff_rdata <= 8'hFF;
			14'd16050: ff_rdata <= 8'hFF;
			14'd16051: ff_rdata <= 8'hFF;
			14'd16052: ff_rdata <= 8'hFF;
			14'd16053: ff_rdata <= 8'hFF;
			14'd16054: ff_rdata <= 8'hFF;
			14'd16055: ff_rdata <= 8'hFF;
			14'd16056: ff_rdata <= 8'hFF;
			14'd16057: ff_rdata <= 8'hFF;
			14'd16058: ff_rdata <= 8'hFF;
			14'd16059: ff_rdata <= 8'hFF;
			14'd16060: ff_rdata <= 8'hFF;
			14'd16061: ff_rdata <= 8'hFF;
			14'd16062: ff_rdata <= 8'hFF;
			14'd16063: ff_rdata <= 8'hFF;
			14'd16064: ff_rdata <= 8'hFF;
			14'd16065: ff_rdata <= 8'hFF;
			14'd16066: ff_rdata <= 8'hFF;
			14'd16067: ff_rdata <= 8'hFF;
			14'd16068: ff_rdata <= 8'hFF;
			14'd16069: ff_rdata <= 8'hFF;
			14'd16070: ff_rdata <= 8'hFF;
			14'd16071: ff_rdata <= 8'hFF;
			14'd16072: ff_rdata <= 8'hFF;
			14'd16073: ff_rdata <= 8'hFF;
			14'd16074: ff_rdata <= 8'hFF;
			14'd16075: ff_rdata <= 8'hFF;
			14'd16076: ff_rdata <= 8'hFF;
			14'd16077: ff_rdata <= 8'hFF;
			14'd16078: ff_rdata <= 8'hFF;
			14'd16079: ff_rdata <= 8'hFF;
			14'd16080: ff_rdata <= 8'hFF;
			14'd16081: ff_rdata <= 8'hFF;
			14'd16082: ff_rdata <= 8'hFF;
			14'd16083: ff_rdata <= 8'hFF;
			14'd16084: ff_rdata <= 8'hFF;
			14'd16085: ff_rdata <= 8'hFF;
			14'd16086: ff_rdata <= 8'hFF;
			14'd16087: ff_rdata <= 8'hFF;
			14'd16088: ff_rdata <= 8'hFF;
			14'd16089: ff_rdata <= 8'hFF;
			14'd16090: ff_rdata <= 8'hFF;
			14'd16091: ff_rdata <= 8'hFF;
			14'd16092: ff_rdata <= 8'hFF;
			14'd16093: ff_rdata <= 8'hFF;
			14'd16094: ff_rdata <= 8'hFF;
			14'd16095: ff_rdata <= 8'hFF;
			14'd16096: ff_rdata <= 8'hFF;
			14'd16097: ff_rdata <= 8'hFF;
			14'd16098: ff_rdata <= 8'hFF;
			14'd16099: ff_rdata <= 8'hFF;
			14'd16100: ff_rdata <= 8'hFF;
			14'd16101: ff_rdata <= 8'hFF;
			14'd16102: ff_rdata <= 8'hFF;
			14'd16103: ff_rdata <= 8'hFF;
			14'd16104: ff_rdata <= 8'hFF;
			14'd16105: ff_rdata <= 8'hFF;
			14'd16106: ff_rdata <= 8'hFF;
			14'd16107: ff_rdata <= 8'hFF;
			14'd16108: ff_rdata <= 8'hFF;
			14'd16109: ff_rdata <= 8'hFF;
			14'd16110: ff_rdata <= 8'hFF;
			14'd16111: ff_rdata <= 8'hFF;
			14'd16112: ff_rdata <= 8'hFF;
			14'd16113: ff_rdata <= 8'hFF;
			14'd16114: ff_rdata <= 8'hFF;
			14'd16115: ff_rdata <= 8'hFF;
			14'd16116: ff_rdata <= 8'hFF;
			14'd16117: ff_rdata <= 8'hFF;
			14'd16118: ff_rdata <= 8'hFF;
			14'd16119: ff_rdata <= 8'hFF;
			14'd16120: ff_rdata <= 8'hFF;
			14'd16121: ff_rdata <= 8'hFF;
			14'd16122: ff_rdata <= 8'hFF;
			14'd16123: ff_rdata <= 8'hFF;
			14'd16124: ff_rdata <= 8'hFF;
			14'd16125: ff_rdata <= 8'hFF;
			14'd16126: ff_rdata <= 8'hFF;
			14'd16127: ff_rdata <= 8'hFF;
			14'd16128: ff_rdata <= 8'hFF;
			14'd16129: ff_rdata <= 8'hFF;
			14'd16130: ff_rdata <= 8'hFF;
			14'd16131: ff_rdata <= 8'hFF;
			14'd16132: ff_rdata <= 8'hFF;
			14'd16133: ff_rdata <= 8'hFF;
			14'd16134: ff_rdata <= 8'hFF;
			14'd16135: ff_rdata <= 8'hFF;
			14'd16136: ff_rdata <= 8'hFF;
			14'd16137: ff_rdata <= 8'hFF;
			14'd16138: ff_rdata <= 8'hFF;
			14'd16139: ff_rdata <= 8'hFF;
			14'd16140: ff_rdata <= 8'hFF;
			14'd16141: ff_rdata <= 8'hFF;
			14'd16142: ff_rdata <= 8'hFF;
			14'd16143: ff_rdata <= 8'hFF;
			14'd16144: ff_rdata <= 8'hFF;
			14'd16145: ff_rdata <= 8'hFF;
			14'd16146: ff_rdata <= 8'hFF;
			14'd16147: ff_rdata <= 8'hFF;
			14'd16148: ff_rdata <= 8'hFF;
			14'd16149: ff_rdata <= 8'hFF;
			14'd16150: ff_rdata <= 8'hFF;
			14'd16151: ff_rdata <= 8'hFF;
			14'd16152: ff_rdata <= 8'hFF;
			14'd16153: ff_rdata <= 8'hFF;
			14'd16154: ff_rdata <= 8'hFF;
			14'd16155: ff_rdata <= 8'hFF;
			14'd16156: ff_rdata <= 8'hFF;
			14'd16157: ff_rdata <= 8'hFF;
			14'd16158: ff_rdata <= 8'hFF;
			14'd16159: ff_rdata <= 8'hFF;
			14'd16160: ff_rdata <= 8'hFF;
			14'd16161: ff_rdata <= 8'hFF;
			14'd16162: ff_rdata <= 8'hFF;
			14'd16163: ff_rdata <= 8'hFF;
			14'd16164: ff_rdata <= 8'hFF;
			14'd16165: ff_rdata <= 8'hFF;
			14'd16166: ff_rdata <= 8'hFF;
			14'd16167: ff_rdata <= 8'hFF;
			14'd16168: ff_rdata <= 8'hFF;
			14'd16169: ff_rdata <= 8'hFF;
			14'd16170: ff_rdata <= 8'hFF;
			14'd16171: ff_rdata <= 8'hFF;
			14'd16172: ff_rdata <= 8'hFF;
			14'd16173: ff_rdata <= 8'hFF;
			14'd16174: ff_rdata <= 8'hFF;
			14'd16175: ff_rdata <= 8'hFF;
			14'd16176: ff_rdata <= 8'hFF;
			14'd16177: ff_rdata <= 8'hFF;
			14'd16178: ff_rdata <= 8'hFF;
			14'd16179: ff_rdata <= 8'hFF;
			14'd16180: ff_rdata <= 8'hFF;
			14'd16181: ff_rdata <= 8'hFF;
			14'd16182: ff_rdata <= 8'hFF;
			14'd16183: ff_rdata <= 8'hFF;
			14'd16184: ff_rdata <= 8'hFF;
			14'd16185: ff_rdata <= 8'hFF;
			14'd16186: ff_rdata <= 8'hFF;
			14'd16187: ff_rdata <= 8'hFF;
			14'd16188: ff_rdata <= 8'hFF;
			14'd16189: ff_rdata <= 8'hFF;
			14'd16190: ff_rdata <= 8'hFF;
			14'd16191: ff_rdata <= 8'hFF;
			14'd16192: ff_rdata <= 8'hFF;
			14'd16193: ff_rdata <= 8'hFF;
			14'd16194: ff_rdata <= 8'hFF;
			14'd16195: ff_rdata <= 8'hFF;
			14'd16196: ff_rdata <= 8'hFF;
			14'd16197: ff_rdata <= 8'hFF;
			14'd16198: ff_rdata <= 8'hFF;
			14'd16199: ff_rdata <= 8'hFF;
			14'd16200: ff_rdata <= 8'hFF;
			14'd16201: ff_rdata <= 8'hFF;
			14'd16202: ff_rdata <= 8'hFF;
			14'd16203: ff_rdata <= 8'hFF;
			14'd16204: ff_rdata <= 8'hFF;
			14'd16205: ff_rdata <= 8'hFF;
			14'd16206: ff_rdata <= 8'hFF;
			14'd16207: ff_rdata <= 8'hFF;
			14'd16208: ff_rdata <= 8'hFF;
			14'd16209: ff_rdata <= 8'hFF;
			14'd16210: ff_rdata <= 8'hFF;
			14'd16211: ff_rdata <= 8'hFF;
			14'd16212: ff_rdata <= 8'hFF;
			14'd16213: ff_rdata <= 8'hFF;
			14'd16214: ff_rdata <= 8'hFF;
			14'd16215: ff_rdata <= 8'hFF;
			14'd16216: ff_rdata <= 8'hFF;
			14'd16217: ff_rdata <= 8'hFF;
			14'd16218: ff_rdata <= 8'hFF;
			14'd16219: ff_rdata <= 8'hFF;
			14'd16220: ff_rdata <= 8'hFF;
			14'd16221: ff_rdata <= 8'hFF;
			14'd16222: ff_rdata <= 8'hFF;
			14'd16223: ff_rdata <= 8'hFF;
			14'd16224: ff_rdata <= 8'hFF;
			14'd16225: ff_rdata <= 8'hFF;
			14'd16226: ff_rdata <= 8'hFF;
			14'd16227: ff_rdata <= 8'hFF;
			14'd16228: ff_rdata <= 8'hFF;
			14'd16229: ff_rdata <= 8'hFF;
			14'd16230: ff_rdata <= 8'hFF;
			14'd16231: ff_rdata <= 8'hFF;
			14'd16232: ff_rdata <= 8'hFF;
			14'd16233: ff_rdata <= 8'hFF;
			14'd16234: ff_rdata <= 8'hFF;
			14'd16235: ff_rdata <= 8'hFF;
			14'd16236: ff_rdata <= 8'hFF;
			14'd16237: ff_rdata <= 8'hFF;
			14'd16238: ff_rdata <= 8'hFF;
			14'd16239: ff_rdata <= 8'hFF;
			14'd16240: ff_rdata <= 8'hFF;
			14'd16241: ff_rdata <= 8'hFF;
			14'd16242: ff_rdata <= 8'hFF;
			14'd16243: ff_rdata <= 8'hFF;
			14'd16244: ff_rdata <= 8'hFF;
			14'd16245: ff_rdata <= 8'hFF;
			14'd16246: ff_rdata <= 8'hFF;
			14'd16247: ff_rdata <= 8'hFF;
			14'd16248: ff_rdata <= 8'hFF;
			14'd16249: ff_rdata <= 8'hFF;
			14'd16250: ff_rdata <= 8'hFF;
			14'd16251: ff_rdata <= 8'hFF;
			14'd16252: ff_rdata <= 8'hFF;
			14'd16253: ff_rdata <= 8'hFF;
			14'd16254: ff_rdata <= 8'hFF;
			14'd16255: ff_rdata <= 8'hFF;
			14'd16256: ff_rdata <= 8'hFF;
			14'd16257: ff_rdata <= 8'hFF;
			14'd16258: ff_rdata <= 8'hFF;
			14'd16259: ff_rdata <= 8'hFF;
			14'd16260: ff_rdata <= 8'hFF;
			14'd16261: ff_rdata <= 8'hFF;
			14'd16262: ff_rdata <= 8'hFF;
			14'd16263: ff_rdata <= 8'hFF;
			14'd16264: ff_rdata <= 8'hFF;
			14'd16265: ff_rdata <= 8'hFF;
			14'd16266: ff_rdata <= 8'hFF;
			14'd16267: ff_rdata <= 8'hFF;
			14'd16268: ff_rdata <= 8'hFF;
			14'd16269: ff_rdata <= 8'hFF;
			14'd16270: ff_rdata <= 8'hFF;
			14'd16271: ff_rdata <= 8'hFF;
			14'd16272: ff_rdata <= 8'hFF;
			14'd16273: ff_rdata <= 8'hFF;
			14'd16274: ff_rdata <= 8'hFF;
			14'd16275: ff_rdata <= 8'hFF;
			14'd16276: ff_rdata <= 8'hFF;
			14'd16277: ff_rdata <= 8'hFF;
			14'd16278: ff_rdata <= 8'hFF;
			14'd16279: ff_rdata <= 8'hFF;
			14'd16280: ff_rdata <= 8'hFF;
			14'd16281: ff_rdata <= 8'hFF;
			14'd16282: ff_rdata <= 8'hFF;
			14'd16283: ff_rdata <= 8'hFF;
			14'd16284: ff_rdata <= 8'hFF;
			14'd16285: ff_rdata <= 8'hFF;
			14'd16286: ff_rdata <= 8'hFF;
			14'd16287: ff_rdata <= 8'hFF;
			14'd16288: ff_rdata <= 8'hFF;
			14'd16289: ff_rdata <= 8'hFF;
			14'd16290: ff_rdata <= 8'hFF;
			14'd16291: ff_rdata <= 8'hFF;
			14'd16292: ff_rdata <= 8'hFF;
			14'd16293: ff_rdata <= 8'hFF;
			14'd16294: ff_rdata <= 8'hFF;
			14'd16295: ff_rdata <= 8'hFF;
			14'd16296: ff_rdata <= 8'hFF;
			14'd16297: ff_rdata <= 8'hFF;
			14'd16298: ff_rdata <= 8'hFF;
			14'd16299: ff_rdata <= 8'hFF;
			14'd16300: ff_rdata <= 8'hFF;
			14'd16301: ff_rdata <= 8'hFF;
			14'd16302: ff_rdata <= 8'hFF;
			14'd16303: ff_rdata <= 8'hFF;
			14'd16304: ff_rdata <= 8'hFF;
			14'd16305: ff_rdata <= 8'hFF;
			14'd16306: ff_rdata <= 8'hFF;
			14'd16307: ff_rdata <= 8'hFF;
			14'd16308: ff_rdata <= 8'hFF;
			14'd16309: ff_rdata <= 8'hFF;
			14'd16310: ff_rdata <= 8'hFF;
			14'd16311: ff_rdata <= 8'hFF;
			14'd16312: ff_rdata <= 8'hFF;
			14'd16313: ff_rdata <= 8'hFF;
			14'd16314: ff_rdata <= 8'hFF;
			14'd16315: ff_rdata <= 8'hFF;
			14'd16316: ff_rdata <= 8'hFF;
			14'd16317: ff_rdata <= 8'hFF;
			14'd16318: ff_rdata <= 8'hFF;
			14'd16319: ff_rdata <= 8'hFF;
			14'd16320: ff_rdata <= 8'hFF;
			14'd16321: ff_rdata <= 8'hFF;
			14'd16322: ff_rdata <= 8'hFF;
			14'd16323: ff_rdata <= 8'hFF;
			14'd16324: ff_rdata <= 8'hFF;
			14'd16325: ff_rdata <= 8'hFF;
			14'd16326: ff_rdata <= 8'hFF;
			14'd16327: ff_rdata <= 8'hFF;
			14'd16328: ff_rdata <= 8'hFF;
			14'd16329: ff_rdata <= 8'hFF;
			14'd16330: ff_rdata <= 8'hFF;
			14'd16331: ff_rdata <= 8'hFF;
			14'd16332: ff_rdata <= 8'hFF;
			14'd16333: ff_rdata <= 8'hFF;
			14'd16334: ff_rdata <= 8'hFF;
			14'd16335: ff_rdata <= 8'hFF;
			14'd16336: ff_rdata <= 8'hFF;
			14'd16337: ff_rdata <= 8'hFF;
			14'd16338: ff_rdata <= 8'hFF;
			14'd16339: ff_rdata <= 8'hFF;
			14'd16340: ff_rdata <= 8'hFF;
			14'd16341: ff_rdata <= 8'hFF;
			14'd16342: ff_rdata <= 8'hFF;
			14'd16343: ff_rdata <= 8'hFF;
			14'd16344: ff_rdata <= 8'hFF;
			14'd16345: ff_rdata <= 8'hFF;
			14'd16346: ff_rdata <= 8'hFF;
			14'd16347: ff_rdata <= 8'hFF;
			14'd16348: ff_rdata <= 8'hFF;
			14'd16349: ff_rdata <= 8'hFF;
			14'd16350: ff_rdata <= 8'hFF;
			14'd16351: ff_rdata <= 8'hFF;
			14'd16352: ff_rdata <= 8'hFF;
			14'd16353: ff_rdata <= 8'hFF;
			14'd16354: ff_rdata <= 8'hFF;
			14'd16355: ff_rdata <= 8'hFF;
			14'd16356: ff_rdata <= 8'hFF;
			14'd16357: ff_rdata <= 8'hFF;
			14'd16358: ff_rdata <= 8'hFF;
			14'd16359: ff_rdata <= 8'hFF;
			14'd16360: ff_rdata <= 8'hFF;
			14'd16361: ff_rdata <= 8'hFF;
			14'd16362: ff_rdata <= 8'hFF;
			14'd16363: ff_rdata <= 8'hFF;
			14'd16364: ff_rdata <= 8'hFF;
			14'd16365: ff_rdata <= 8'hC3;
			14'd16366: ff_rdata <= 8'h03;
			14'd16367: ff_rdata <= 8'h50;
			14'd16368: ff_rdata <= 8'hFF;
			14'd16369: ff_rdata <= 8'hFF;
			14'd16370: ff_rdata <= 8'hFF;
			14'd16371: ff_rdata <= 8'hFF;
			14'd16372: ff_rdata <= 8'hFF;
			14'd16373: ff_rdata <= 8'hFF;
			14'd16374: ff_rdata <= 8'h00;
			14'd16375: ff_rdata <= 8'h00;
			14'd16376: ff_rdata <= 8'hFF;
			14'd16377: ff_rdata <= 8'hFF;
			14'd16378: ff_rdata <= 8'hFF;
			14'd16379: ff_rdata <= 8'hFF;
			14'd16380: ff_rdata <= 8'hFF;
			14'd16381: ff_rdata <= 8'hFF;
			14'd16382: ff_rdata <= 8'hFF;
			14'd16383: ff_rdata <= 8'hFF;
			default: ff_rdata <= 8'd0;
			endcase
			ff_rdata_en <= 1'b1;
		end
		else begin
			ff_rdata <= 8'd0;
			ff_rdata_en <= 1'b0;
		end
	end

	assign rdata	= ff_rdata;
	assign rdata_en	= ff_rdata_en;
endmodule
