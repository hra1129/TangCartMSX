reg [7:0] ff_ram [0:16383];
initial begin
    ff_ram[0] = 8'h00;
    ff_ram[1] = 8'h00;
    ff_ram[2] = 8'h00;
    ff_ram[3] = 8'h00;
    ff_ram[4] = 8'h00;
    ff_ram[5] = 8'h00;
    ff_ram[6] = 8'h00;
    ff_ram[7] = 8'h00;
    ff_ram[8] = 8'h7E;
    ff_ram[9] = 8'h42;
    ff_ram[10] = 8'h7E;
    ff_ram[11] = 8'h42;
    ff_ram[12] = 8'h7E;
    ff_ram[13] = 8'h42;
    ff_ram[14] = 8'h82;
    ff_ram[15] = 8'h00;
    ff_ram[16] = 8'h10;
    ff_ram[17] = 8'h92;
    ff_ram[18] = 8'h54;
    ff_ram[19] = 8'h10;
    ff_ram[20] = 8'h28;
    ff_ram[21] = 8'h44;
    ff_ram[22] = 8'h82;
    ff_ram[23] = 8'h00;
    ff_ram[24] = 8'h12;
    ff_ram[25] = 8'h14;
    ff_ram[26] = 8'hF8;
    ff_ram[27] = 8'h14;
    ff_ram[28] = 8'h34;
    ff_ram[29] = 8'h52;
    ff_ram[30] = 8'h92;
    ff_ram[31] = 8'h00;
    ff_ram[32] = 8'h10;
    ff_ram[33] = 8'h10;
    ff_ram[34] = 8'hFE;
    ff_ram[35] = 8'h10;
    ff_ram[36] = 8'h38;
    ff_ram[37] = 8'h54;
    ff_ram[38] = 8'h92;
    ff_ram[39] = 8'h00;
    ff_ram[40] = 8'h10;
    ff_ram[41] = 8'h28;
    ff_ram[42] = 8'h7C;
    ff_ram[43] = 8'h92;
    ff_ram[44] = 8'h38;
    ff_ram[45] = 8'h54;
    ff_ram[46] = 8'hFE;
    ff_ram[47] = 8'h00;
    ff_ram[48] = 8'h10;
    ff_ram[49] = 8'h10;
    ff_ram[50] = 8'h10;
    ff_ram[51] = 8'h7C;
    ff_ram[52] = 8'h10;
    ff_ram[53] = 8'h10;
    ff_ram[54] = 8'hFE;
    ff_ram[55] = 8'h00;
    ff_ram[56] = 8'h7E;
    ff_ram[57] = 8'h42;
    ff_ram[58] = 8'h42;
    ff_ram[59] = 8'h7E;
    ff_ram[60] = 8'h42;
    ff_ram[61] = 8'h42;
    ff_ram[62] = 8'h7E;
    ff_ram[63] = 8'h00;
    ff_ram[64] = 8'h40;
    ff_ram[65] = 8'h7E;
    ff_ram[66] = 8'h48;
    ff_ram[67] = 8'h3C;
    ff_ram[68] = 8'h28;
    ff_ram[69] = 8'h7E;
    ff_ram[70] = 8'h08;
    ff_ram[71] = 8'h00;
    ff_ram[72] = 8'hFE;
    ff_ram[73] = 8'h92;
    ff_ram[74] = 8'h92;
    ff_ram[75] = 8'hFE;
    ff_ram[76] = 8'h82;
    ff_ram[77] = 8'h82;
    ff_ram[78] = 8'h86;
    ff_ram[79] = 8'h00;
    ff_ram[80] = 8'h04;
    ff_ram[81] = 8'hEE;
    ff_ram[82] = 8'hA4;
    ff_ram[83] = 8'hEF;
    ff_ram[84] = 8'hA2;
    ff_ram[85] = 8'hEA;
    ff_ram[86] = 8'h06;
    ff_ram[87] = 8'h00;
    ff_ram[88] = 8'h28;
    ff_ram[89] = 8'h44;
    ff_ram[90] = 8'h82;
    ff_ram[91] = 8'h3C;
    ff_ram[92] = 8'h14;
    ff_ram[93] = 8'h24;
    ff_ram[94] = 8'h4C;
    ff_ram[95] = 8'h00;
    ff_ram[96] = 8'h28;
    ff_ram[97] = 8'hC8;
    ff_ram[98] = 8'h5C;
    ff_ram[99] = 8'hEA;
    ff_ram[100] = 8'h6C;
    ff_ram[101] = 8'hC8;
    ff_ram[102] = 8'h50;
    ff_ram[103] = 8'h00;
    ff_ram[104] = 8'h7C;
    ff_ram[105] = 8'h20;
    ff_ram[106] = 8'h7C;
    ff_ram[107] = 8'h44;
    ff_ram[108] = 8'h7C;
    ff_ram[109] = 8'h44;
    ff_ram[110] = 8'h7C;
    ff_ram[111] = 8'h00;
    ff_ram[112] = 8'h0C;
    ff_ram[113] = 8'h70;
    ff_ram[114] = 8'h10;
    ff_ram[115] = 8'hFE;
    ff_ram[116] = 8'h10;
    ff_ram[117] = 8'h10;
    ff_ram[118] = 8'h10;
    ff_ram[119] = 8'h00;
    ff_ram[120] = 8'h7E;
    ff_ram[121] = 8'h10;
    ff_ram[122] = 8'h1E;
    ff_ram[123] = 8'h12;
    ff_ram[124] = 8'h22;
    ff_ram[125] = 8'h44;
    ff_ram[126] = 8'h08;
    ff_ram[127] = 8'h00;
    ff_ram[128] = 8'h00;
    ff_ram[129] = 8'h7C;
    ff_ram[130] = 8'h28;
    ff_ram[131] = 8'h28;
    ff_ram[132] = 8'h28;
    ff_ram[133] = 8'h4E;
    ff_ram[134] = 8'h00;
    ff_ram[135] = 8'h00;
    ff_ram[136] = 8'h10;
    ff_ram[137] = 8'h10;
    ff_ram[138] = 8'h10;
    ff_ram[139] = 8'hFF;
    ff_ram[140] = 8'h00;
    ff_ram[141] = 8'h00;
    ff_ram[142] = 8'h00;
    ff_ram[143] = 8'h00;
    ff_ram[144] = 8'h00;
    ff_ram[145] = 8'h00;
    ff_ram[146] = 8'h00;
    ff_ram[147] = 8'hFF;
    ff_ram[148] = 8'h10;
    ff_ram[149] = 8'h10;
    ff_ram[150] = 8'h10;
    ff_ram[151] = 8'h10;
    ff_ram[152] = 8'h10;
    ff_ram[153] = 8'h10;
    ff_ram[154] = 8'h10;
    ff_ram[155] = 8'hF0;
    ff_ram[156] = 8'h10;
    ff_ram[157] = 8'h10;
    ff_ram[158] = 8'h10;
    ff_ram[159] = 8'h10;
    ff_ram[160] = 8'h10;
    ff_ram[161] = 8'h10;
    ff_ram[162] = 8'h10;
    ff_ram[163] = 8'h1F;
    ff_ram[164] = 8'h10;
    ff_ram[165] = 8'h10;
    ff_ram[166] = 8'h10;
    ff_ram[167] = 8'h10;
    ff_ram[168] = 8'h10;
    ff_ram[169] = 8'h10;
    ff_ram[170] = 8'h10;
    ff_ram[171] = 8'hFF;
    ff_ram[172] = 8'h10;
    ff_ram[173] = 8'h10;
    ff_ram[174] = 8'h10;
    ff_ram[175] = 8'h10;
    ff_ram[176] = 8'h10;
    ff_ram[177] = 8'h10;
    ff_ram[178] = 8'h10;
    ff_ram[179] = 8'h10;
    ff_ram[180] = 8'h10;
    ff_ram[181] = 8'h10;
    ff_ram[182] = 8'h10;
    ff_ram[183] = 8'h10;
    ff_ram[184] = 8'h00;
    ff_ram[185] = 8'h00;
    ff_ram[186] = 8'h00;
    ff_ram[187] = 8'hFF;
    ff_ram[188] = 8'h00;
    ff_ram[189] = 8'h00;
    ff_ram[190] = 8'h00;
    ff_ram[191] = 8'h00;
    ff_ram[192] = 8'h00;
    ff_ram[193] = 8'h00;
    ff_ram[194] = 8'h00;
    ff_ram[195] = 8'h1F;
    ff_ram[196] = 8'h10;
    ff_ram[197] = 8'h10;
    ff_ram[198] = 8'h10;
    ff_ram[199] = 8'h10;
    ff_ram[200] = 8'h00;
    ff_ram[201] = 8'h00;
    ff_ram[202] = 8'h00;
    ff_ram[203] = 8'hF0;
    ff_ram[204] = 8'h10;
    ff_ram[205] = 8'h10;
    ff_ram[206] = 8'h10;
    ff_ram[207] = 8'h10;
    ff_ram[208] = 8'h10;
    ff_ram[209] = 8'h10;
    ff_ram[210] = 8'h10;
    ff_ram[211] = 8'h1F;
    ff_ram[212] = 8'h00;
    ff_ram[213] = 8'h00;
    ff_ram[214] = 8'h00;
    ff_ram[215] = 8'h00;
    ff_ram[216] = 8'h10;
    ff_ram[217] = 8'h10;
    ff_ram[218] = 8'h10;
    ff_ram[219] = 8'hF0;
    ff_ram[220] = 8'h00;
    ff_ram[221] = 8'h00;
    ff_ram[222] = 8'h00;
    ff_ram[223] = 8'h00;
    ff_ram[224] = 8'h81;
    ff_ram[225] = 8'h42;
    ff_ram[226] = 8'h24;
    ff_ram[227] = 8'h18;
    ff_ram[228] = 8'h18;
    ff_ram[229] = 8'h24;
    ff_ram[230] = 8'h42;
    ff_ram[231] = 8'h81;
    ff_ram[232] = 8'h10;
    ff_ram[233] = 8'h7C;
    ff_ram[234] = 8'h10;
    ff_ram[235] = 8'h10;
    ff_ram[236] = 8'h28;
    ff_ram[237] = 8'h44;
    ff_ram[238] = 8'h82;
    ff_ram[239] = 8'h00;
    ff_ram[240] = 8'h10;
    ff_ram[241] = 8'h10;
    ff_ram[242] = 8'hFE;
    ff_ram[243] = 8'h92;
    ff_ram[244] = 8'hFE;
    ff_ram[245] = 8'h10;
    ff_ram[246] = 8'h10;
    ff_ram[247] = 8'h00;
    ff_ram[248] = 8'h10;
    ff_ram[249] = 8'h10;
    ff_ram[250] = 8'h54;
    ff_ram[251] = 8'h54;
    ff_ram[252] = 8'h92;
    ff_ram[253] = 8'h10;
    ff_ram[254] = 8'h30;
    ff_ram[255] = 8'h00;
    ff_ram[256] = 8'h00;
    ff_ram[257] = 8'h00;
    ff_ram[258] = 8'h00;
    ff_ram[259] = 8'h00;
    ff_ram[260] = 8'h00;
    ff_ram[261] = 8'h00;
    ff_ram[262] = 8'h00;
    ff_ram[263] = 8'h00;
    ff_ram[264] = 8'h20;
    ff_ram[265] = 8'h20;
    ff_ram[266] = 8'h20;
    ff_ram[267] = 8'h20;
    ff_ram[268] = 8'h00;
    ff_ram[269] = 8'h00;
    ff_ram[270] = 8'h20;
    ff_ram[271] = 8'h00;
    ff_ram[272] = 8'h50;
    ff_ram[273] = 8'h50;
    ff_ram[274] = 8'h50;
    ff_ram[275] = 8'h00;
    ff_ram[276] = 8'h00;
    ff_ram[277] = 8'h00;
    ff_ram[278] = 8'h00;
    ff_ram[279] = 8'h00;
    ff_ram[280] = 8'h50;
    ff_ram[281] = 8'h50;
    ff_ram[282] = 8'hF8;
    ff_ram[283] = 8'h50;
    ff_ram[284] = 8'hF8;
    ff_ram[285] = 8'h50;
    ff_ram[286] = 8'h50;
    ff_ram[287] = 8'h00;
    ff_ram[288] = 8'h20;
    ff_ram[289] = 8'h78;
    ff_ram[290] = 8'hA0;
    ff_ram[291] = 8'h70;
    ff_ram[292] = 8'h28;
    ff_ram[293] = 8'hF0;
    ff_ram[294] = 8'h20;
    ff_ram[295] = 8'h00;
    ff_ram[296] = 8'hC0;
    ff_ram[297] = 8'hC8;
    ff_ram[298] = 8'h10;
    ff_ram[299] = 8'h20;
    ff_ram[300] = 8'h40;
    ff_ram[301] = 8'h98;
    ff_ram[302] = 8'h18;
    ff_ram[303] = 8'h00;
    ff_ram[304] = 8'h40;
    ff_ram[305] = 8'hA0;
    ff_ram[306] = 8'h40;
    ff_ram[307] = 8'hA8;
    ff_ram[308] = 8'h90;
    ff_ram[309] = 8'h98;
    ff_ram[310] = 8'h60;
    ff_ram[311] = 8'h00;
    ff_ram[312] = 8'h10;
    ff_ram[313] = 8'h20;
    ff_ram[314] = 8'h40;
    ff_ram[315] = 8'h00;
    ff_ram[316] = 8'h00;
    ff_ram[317] = 8'h00;
    ff_ram[318] = 8'h00;
    ff_ram[319] = 8'h00;
    ff_ram[320] = 8'h10;
    ff_ram[321] = 8'h20;
    ff_ram[322] = 8'h40;
    ff_ram[323] = 8'h40;
    ff_ram[324] = 8'h40;
    ff_ram[325] = 8'h20;
    ff_ram[326] = 8'h10;
    ff_ram[327] = 8'h00;
    ff_ram[328] = 8'h40;
    ff_ram[329] = 8'h20;
    ff_ram[330] = 8'h10;
    ff_ram[331] = 8'h10;
    ff_ram[332] = 8'h10;
    ff_ram[333] = 8'h20;
    ff_ram[334] = 8'h40;
    ff_ram[335] = 8'h00;
    ff_ram[336] = 8'h20;
    ff_ram[337] = 8'hA8;
    ff_ram[338] = 8'h70;
    ff_ram[339] = 8'h20;
    ff_ram[340] = 8'h70;
    ff_ram[341] = 8'hA8;
    ff_ram[342] = 8'h20;
    ff_ram[343] = 8'h00;
    ff_ram[344] = 8'h00;
    ff_ram[345] = 8'h20;
    ff_ram[346] = 8'h20;
    ff_ram[347] = 8'hF8;
    ff_ram[348] = 8'h20;
    ff_ram[349] = 8'h20;
    ff_ram[350] = 8'h00;
    ff_ram[351] = 8'h00;
    ff_ram[352] = 8'h00;
    ff_ram[353] = 8'h00;
    ff_ram[354] = 8'h00;
    ff_ram[355] = 8'h00;
    ff_ram[356] = 8'h00;
    ff_ram[357] = 8'h20;
    ff_ram[358] = 8'h20;
    ff_ram[359] = 8'h40;
    ff_ram[360] = 8'h00;
    ff_ram[361] = 8'h00;
    ff_ram[362] = 8'h00;
    ff_ram[363] = 8'h78;
    ff_ram[364] = 8'h00;
    ff_ram[365] = 8'h00;
    ff_ram[366] = 8'h00;
    ff_ram[367] = 8'h00;
    ff_ram[368] = 8'h00;
    ff_ram[369] = 8'h00;
    ff_ram[370] = 8'h00;
    ff_ram[371] = 8'h00;
    ff_ram[372] = 8'h00;
    ff_ram[373] = 8'h60;
    ff_ram[374] = 8'h60;
    ff_ram[375] = 8'h00;
    ff_ram[376] = 8'h00;
    ff_ram[377] = 8'h00;
    ff_ram[378] = 8'h08;
    ff_ram[379] = 8'h10;
    ff_ram[380] = 8'h20;
    ff_ram[381] = 8'h40;
    ff_ram[382] = 8'h80;
    ff_ram[383] = 8'h00;
    ff_ram[384] = 8'h70;
    ff_ram[385] = 8'h88;
    ff_ram[386] = 8'h98;
    ff_ram[387] = 8'hA8;
    ff_ram[388] = 8'hC8;
    ff_ram[389] = 8'h88;
    ff_ram[390] = 8'h70;
    ff_ram[391] = 8'h00;
    ff_ram[392] = 8'h20;
    ff_ram[393] = 8'h60;
    ff_ram[394] = 8'hA0;
    ff_ram[395] = 8'h20;
    ff_ram[396] = 8'h20;
    ff_ram[397] = 8'h20;
    ff_ram[398] = 8'hF8;
    ff_ram[399] = 8'h00;
    ff_ram[400] = 8'h70;
    ff_ram[401] = 8'h88;
    ff_ram[402] = 8'h08;
    ff_ram[403] = 8'h10;
    ff_ram[404] = 8'h60;
    ff_ram[405] = 8'h80;
    ff_ram[406] = 8'hF8;
    ff_ram[407] = 8'h00;
    ff_ram[408] = 8'h70;
    ff_ram[409] = 8'h88;
    ff_ram[410] = 8'h08;
    ff_ram[411] = 8'h30;
    ff_ram[412] = 8'h08;
    ff_ram[413] = 8'h88;
    ff_ram[414] = 8'h70;
    ff_ram[415] = 8'h00;
    ff_ram[416] = 8'h10;
    ff_ram[417] = 8'h30;
    ff_ram[418] = 8'h50;
    ff_ram[419] = 8'h90;
    ff_ram[420] = 8'hF8;
    ff_ram[421] = 8'h10;
    ff_ram[422] = 8'h10;
    ff_ram[423] = 8'h00;
    ff_ram[424] = 8'hF8;
    ff_ram[425] = 8'h80;
    ff_ram[426] = 8'hE0;
    ff_ram[427] = 8'h10;
    ff_ram[428] = 8'h08;
    ff_ram[429] = 8'h10;
    ff_ram[430] = 8'hE0;
    ff_ram[431] = 8'h00;
    ff_ram[432] = 8'h30;
    ff_ram[433] = 8'h40;
    ff_ram[434] = 8'h80;
    ff_ram[435] = 8'hF0;
    ff_ram[436] = 8'h88;
    ff_ram[437] = 8'h88;
    ff_ram[438] = 8'h70;
    ff_ram[439] = 8'h00;
    ff_ram[440] = 8'hF8;
    ff_ram[441] = 8'h88;
    ff_ram[442] = 8'h10;
    ff_ram[443] = 8'h20;
    ff_ram[444] = 8'h20;
    ff_ram[445] = 8'h20;
    ff_ram[446] = 8'h20;
    ff_ram[447] = 8'h00;
    ff_ram[448] = 8'h70;
    ff_ram[449] = 8'h88;
    ff_ram[450] = 8'h88;
    ff_ram[451] = 8'h70;
    ff_ram[452] = 8'h88;
    ff_ram[453] = 8'h88;
    ff_ram[454] = 8'h70;
    ff_ram[455] = 8'h00;
    ff_ram[456] = 8'h70;
    ff_ram[457] = 8'h88;
    ff_ram[458] = 8'h88;
    ff_ram[459] = 8'h78;
    ff_ram[460] = 8'h08;
    ff_ram[461] = 8'h10;
    ff_ram[462] = 8'h60;
    ff_ram[463] = 8'h00;
    ff_ram[464] = 8'h00;
    ff_ram[465] = 8'h00;
    ff_ram[466] = 8'h20;
    ff_ram[467] = 8'h00;
    ff_ram[468] = 8'h00;
    ff_ram[469] = 8'h20;
    ff_ram[470] = 8'h00;
    ff_ram[471] = 8'h00;
    ff_ram[472] = 8'h00;
    ff_ram[473] = 8'h00;
    ff_ram[474] = 8'h20;
    ff_ram[475] = 8'h00;
    ff_ram[476] = 8'h00;
    ff_ram[477] = 8'h20;
    ff_ram[478] = 8'h20;
    ff_ram[479] = 8'h40;
    ff_ram[480] = 8'h18;
    ff_ram[481] = 8'h30;
    ff_ram[482] = 8'h60;
    ff_ram[483] = 8'hC0;
    ff_ram[484] = 8'h60;
    ff_ram[485] = 8'h30;
    ff_ram[486] = 8'h18;
    ff_ram[487] = 8'h00;
    ff_ram[488] = 8'h00;
    ff_ram[489] = 8'h00;
    ff_ram[490] = 8'hF8;
    ff_ram[491] = 8'h00;
    ff_ram[492] = 8'hF8;
    ff_ram[493] = 8'h00;
    ff_ram[494] = 8'h00;
    ff_ram[495] = 8'h00;
    ff_ram[496] = 8'hC0;
    ff_ram[497] = 8'h60;
    ff_ram[498] = 8'h30;
    ff_ram[499] = 8'h18;
    ff_ram[500] = 8'h30;
    ff_ram[501] = 8'h60;
    ff_ram[502] = 8'hC0;
    ff_ram[503] = 8'h00;
    ff_ram[504] = 8'h70;
    ff_ram[505] = 8'h88;
    ff_ram[506] = 8'h08;
    ff_ram[507] = 8'h10;
    ff_ram[508] = 8'h20;
    ff_ram[509] = 8'h00;
    ff_ram[510] = 8'h20;
    ff_ram[511] = 8'h00;
    ff_ram[512] = 8'h70;
    ff_ram[513] = 8'h88;
    ff_ram[514] = 8'h08;
    ff_ram[515] = 8'h68;
    ff_ram[516] = 8'hA8;
    ff_ram[517] = 8'hA8;
    ff_ram[518] = 8'h70;
    ff_ram[519] = 8'h00;
    ff_ram[520] = 8'h20;
    ff_ram[521] = 8'h50;
    ff_ram[522] = 8'h88;
    ff_ram[523] = 8'h88;
    ff_ram[524] = 8'hF8;
    ff_ram[525] = 8'h88;
    ff_ram[526] = 8'h88;
    ff_ram[527] = 8'h00;
    ff_ram[528] = 8'hF0;
    ff_ram[529] = 8'h48;
    ff_ram[530] = 8'h48;
    ff_ram[531] = 8'h70;
    ff_ram[532] = 8'h48;
    ff_ram[533] = 8'h48;
    ff_ram[534] = 8'hF0;
    ff_ram[535] = 8'h00;
    ff_ram[536] = 8'h30;
    ff_ram[537] = 8'h48;
    ff_ram[538] = 8'h80;
    ff_ram[539] = 8'h80;
    ff_ram[540] = 8'h80;
    ff_ram[541] = 8'h48;
    ff_ram[542] = 8'h30;
    ff_ram[543] = 8'h00;
    ff_ram[544] = 8'hE0;
    ff_ram[545] = 8'h50;
    ff_ram[546] = 8'h48;
    ff_ram[547] = 8'h48;
    ff_ram[548] = 8'h48;
    ff_ram[549] = 8'h50;
    ff_ram[550] = 8'hE0;
    ff_ram[551] = 8'h00;
    ff_ram[552] = 8'hF8;
    ff_ram[553] = 8'h80;
    ff_ram[554] = 8'h80;
    ff_ram[555] = 8'hF0;
    ff_ram[556] = 8'h80;
    ff_ram[557] = 8'h80;
    ff_ram[558] = 8'hF8;
    ff_ram[559] = 8'h00;
    ff_ram[560] = 8'hF8;
    ff_ram[561] = 8'h80;
    ff_ram[562] = 8'h80;
    ff_ram[563] = 8'hF0;
    ff_ram[564] = 8'h80;
    ff_ram[565] = 8'h80;
    ff_ram[566] = 8'h80;
    ff_ram[567] = 8'h00;
    ff_ram[568] = 8'h70;
    ff_ram[569] = 8'h88;
    ff_ram[570] = 8'h80;
    ff_ram[571] = 8'hB8;
    ff_ram[572] = 8'h88;
    ff_ram[573] = 8'h88;
    ff_ram[574] = 8'h70;
    ff_ram[575] = 8'h00;
    ff_ram[576] = 8'h88;
    ff_ram[577] = 8'h88;
    ff_ram[578] = 8'h88;
    ff_ram[579] = 8'hF8;
    ff_ram[580] = 8'h88;
    ff_ram[581] = 8'h88;
    ff_ram[582] = 8'h88;
    ff_ram[583] = 8'h00;
    ff_ram[584] = 8'h70;
    ff_ram[585] = 8'h20;
    ff_ram[586] = 8'h20;
    ff_ram[587] = 8'h20;
    ff_ram[588] = 8'h20;
    ff_ram[589] = 8'h20;
    ff_ram[590] = 8'h70;
    ff_ram[591] = 8'h00;
    ff_ram[592] = 8'h38;
    ff_ram[593] = 8'h10;
    ff_ram[594] = 8'h10;
    ff_ram[595] = 8'h10;
    ff_ram[596] = 8'h90;
    ff_ram[597] = 8'h90;
    ff_ram[598] = 8'h60;
    ff_ram[599] = 8'h00;
    ff_ram[600] = 8'h88;
    ff_ram[601] = 8'h90;
    ff_ram[602] = 8'hA0;
    ff_ram[603] = 8'hC0;
    ff_ram[604] = 8'hA0;
    ff_ram[605] = 8'h90;
    ff_ram[606] = 8'h88;
    ff_ram[607] = 8'h00;
    ff_ram[608] = 8'h80;
    ff_ram[609] = 8'h80;
    ff_ram[610] = 8'h80;
    ff_ram[611] = 8'h80;
    ff_ram[612] = 8'h80;
    ff_ram[613] = 8'h80;
    ff_ram[614] = 8'hF8;
    ff_ram[615] = 8'h00;
    ff_ram[616] = 8'h88;
    ff_ram[617] = 8'hD8;
    ff_ram[618] = 8'hA8;
    ff_ram[619] = 8'hA8;
    ff_ram[620] = 8'h88;
    ff_ram[621] = 8'h88;
    ff_ram[622] = 8'h88;
    ff_ram[623] = 8'h00;
    ff_ram[624] = 8'h88;
    ff_ram[625] = 8'hC8;
    ff_ram[626] = 8'hC8;
    ff_ram[627] = 8'hA8;
    ff_ram[628] = 8'h98;
    ff_ram[629] = 8'h98;
    ff_ram[630] = 8'h88;
    ff_ram[631] = 8'h00;
    ff_ram[632] = 8'h70;
    ff_ram[633] = 8'h88;
    ff_ram[634] = 8'h88;
    ff_ram[635] = 8'h88;
    ff_ram[636] = 8'h88;
    ff_ram[637] = 8'h88;
    ff_ram[638] = 8'h70;
    ff_ram[639] = 8'h00;
    ff_ram[640] = 8'hF0;
    ff_ram[641] = 8'h88;
    ff_ram[642] = 8'h88;
    ff_ram[643] = 8'hF0;
    ff_ram[644] = 8'h80;
    ff_ram[645] = 8'h80;
    ff_ram[646] = 8'h80;
    ff_ram[647] = 8'h00;
    ff_ram[648] = 8'h70;
    ff_ram[649] = 8'h88;
    ff_ram[650] = 8'h88;
    ff_ram[651] = 8'h88;
    ff_ram[652] = 8'hA8;
    ff_ram[653] = 8'h90;
    ff_ram[654] = 8'h68;
    ff_ram[655] = 8'h00;
    ff_ram[656] = 8'hF0;
    ff_ram[657] = 8'h88;
    ff_ram[658] = 8'h88;
    ff_ram[659] = 8'hF0;
    ff_ram[660] = 8'hA0;
    ff_ram[661] = 8'h90;
    ff_ram[662] = 8'h88;
    ff_ram[663] = 8'h00;
    ff_ram[664] = 8'h70;
    ff_ram[665] = 8'h88;
    ff_ram[666] = 8'h80;
    ff_ram[667] = 8'h70;
    ff_ram[668] = 8'h08;
    ff_ram[669] = 8'h88;
    ff_ram[670] = 8'h70;
    ff_ram[671] = 8'h00;
    ff_ram[672] = 8'hF8;
    ff_ram[673] = 8'h20;
    ff_ram[674] = 8'h20;
    ff_ram[675] = 8'h20;
    ff_ram[676] = 8'h20;
    ff_ram[677] = 8'h20;
    ff_ram[678] = 8'h20;
    ff_ram[679] = 8'h00;
    ff_ram[680] = 8'h88;
    ff_ram[681] = 8'h88;
    ff_ram[682] = 8'h88;
    ff_ram[683] = 8'h88;
    ff_ram[684] = 8'h88;
    ff_ram[685] = 8'h88;
    ff_ram[686] = 8'h70;
    ff_ram[687] = 8'h00;
    ff_ram[688] = 8'h88;
    ff_ram[689] = 8'h88;
    ff_ram[690] = 8'h88;
    ff_ram[691] = 8'h88;
    ff_ram[692] = 8'h50;
    ff_ram[693] = 8'h50;
    ff_ram[694] = 8'h20;
    ff_ram[695] = 8'h00;
    ff_ram[696] = 8'h88;
    ff_ram[697] = 8'h88;
    ff_ram[698] = 8'h88;
    ff_ram[699] = 8'hA8;
    ff_ram[700] = 8'hA8;
    ff_ram[701] = 8'hD8;
    ff_ram[702] = 8'h88;
    ff_ram[703] = 8'h00;
    ff_ram[704] = 8'h88;
    ff_ram[705] = 8'h88;
    ff_ram[706] = 8'h50;
    ff_ram[707] = 8'h20;
    ff_ram[708] = 8'h50;
    ff_ram[709] = 8'h88;
    ff_ram[710] = 8'h88;
    ff_ram[711] = 8'h00;
    ff_ram[712] = 8'h88;
    ff_ram[713] = 8'h88;
    ff_ram[714] = 8'h88;
    ff_ram[715] = 8'h70;
    ff_ram[716] = 8'h20;
    ff_ram[717] = 8'h20;
    ff_ram[718] = 8'h20;
    ff_ram[719] = 8'h00;
    ff_ram[720] = 8'hF8;
    ff_ram[721] = 8'h08;
    ff_ram[722] = 8'h10;
    ff_ram[723] = 8'h20;
    ff_ram[724] = 8'h40;
    ff_ram[725] = 8'h80;
    ff_ram[726] = 8'hF8;
    ff_ram[727] = 8'h00;
    ff_ram[728] = 8'h70;
    ff_ram[729] = 8'h40;
    ff_ram[730] = 8'h40;
    ff_ram[731] = 8'h40;
    ff_ram[732] = 8'h40;
    ff_ram[733] = 8'h40;
    ff_ram[734] = 8'h70;
    ff_ram[735] = 8'h00;
    ff_ram[736] = 8'h88;
    ff_ram[737] = 8'h50;
    ff_ram[738] = 8'h20;
    ff_ram[739] = 8'h70;
    ff_ram[740] = 8'h20;
    ff_ram[741] = 8'h70;
    ff_ram[742] = 8'h20;
    ff_ram[743] = 8'h00;
    ff_ram[744] = 8'h70;
    ff_ram[745] = 8'h10;
    ff_ram[746] = 8'h10;
    ff_ram[747] = 8'h10;
    ff_ram[748] = 8'h10;
    ff_ram[749] = 8'h10;
    ff_ram[750] = 8'h70;
    ff_ram[751] = 8'h00;
    ff_ram[752] = 8'h20;
    ff_ram[753] = 8'h50;
    ff_ram[754] = 8'h88;
    ff_ram[755] = 8'h00;
    ff_ram[756] = 8'h00;
    ff_ram[757] = 8'h00;
    ff_ram[758] = 8'h00;
    ff_ram[759] = 8'h00;
    ff_ram[760] = 8'h00;
    ff_ram[761] = 8'h00;
    ff_ram[762] = 8'h00;
    ff_ram[763] = 8'h00;
    ff_ram[764] = 8'h00;
    ff_ram[765] = 8'h00;
    ff_ram[766] = 8'hF8;
    ff_ram[767] = 8'h00;
    ff_ram[768] = 8'h40;
    ff_ram[769] = 8'h20;
    ff_ram[770] = 8'h10;
    ff_ram[771] = 8'h00;
    ff_ram[772] = 8'h00;
    ff_ram[773] = 8'h00;
    ff_ram[774] = 8'h00;
    ff_ram[775] = 8'h00;
    ff_ram[776] = 8'h00;
    ff_ram[777] = 8'h00;
    ff_ram[778] = 8'h70;
    ff_ram[779] = 8'h08;
    ff_ram[780] = 8'h78;
    ff_ram[781] = 8'h88;
    ff_ram[782] = 8'h78;
    ff_ram[783] = 8'h00;
    ff_ram[784] = 8'h80;
    ff_ram[785] = 8'h80;
    ff_ram[786] = 8'hB0;
    ff_ram[787] = 8'hC8;
    ff_ram[788] = 8'h88;
    ff_ram[789] = 8'hC8;
    ff_ram[790] = 8'hB0;
    ff_ram[791] = 8'h00;
    ff_ram[792] = 8'h00;
    ff_ram[793] = 8'h00;
    ff_ram[794] = 8'h70;
    ff_ram[795] = 8'h88;
    ff_ram[796] = 8'h80;
    ff_ram[797] = 8'h88;
    ff_ram[798] = 8'h70;
    ff_ram[799] = 8'h00;
    ff_ram[800] = 8'h08;
    ff_ram[801] = 8'h08;
    ff_ram[802] = 8'h68;
    ff_ram[803] = 8'h98;
    ff_ram[804] = 8'h88;
    ff_ram[805] = 8'h98;
    ff_ram[806] = 8'h68;
    ff_ram[807] = 8'h00;
    ff_ram[808] = 8'h00;
    ff_ram[809] = 8'h00;
    ff_ram[810] = 8'h70;
    ff_ram[811] = 8'h88;
    ff_ram[812] = 8'hF8;
    ff_ram[813] = 8'h80;
    ff_ram[814] = 8'h70;
    ff_ram[815] = 8'h00;
    ff_ram[816] = 8'h10;
    ff_ram[817] = 8'h28;
    ff_ram[818] = 8'h20;
    ff_ram[819] = 8'hF8;
    ff_ram[820] = 8'h20;
    ff_ram[821] = 8'h20;
    ff_ram[822] = 8'h20;
    ff_ram[823] = 8'h00;
    ff_ram[824] = 8'h00;
    ff_ram[825] = 8'h00;
    ff_ram[826] = 8'h68;
    ff_ram[827] = 8'h98;
    ff_ram[828] = 8'h98;
    ff_ram[829] = 8'h68;
    ff_ram[830] = 8'h08;
    ff_ram[831] = 8'h70;
    ff_ram[832] = 8'h80;
    ff_ram[833] = 8'h80;
    ff_ram[834] = 8'hF0;
    ff_ram[835] = 8'h88;
    ff_ram[836] = 8'h88;
    ff_ram[837] = 8'h88;
    ff_ram[838] = 8'h88;
    ff_ram[839] = 8'h00;
    ff_ram[840] = 8'h20;
    ff_ram[841] = 8'h00;
    ff_ram[842] = 8'h60;
    ff_ram[843] = 8'h20;
    ff_ram[844] = 8'h20;
    ff_ram[845] = 8'h20;
    ff_ram[846] = 8'h70;
    ff_ram[847] = 8'h00;
    ff_ram[848] = 8'h10;
    ff_ram[849] = 8'h00;
    ff_ram[850] = 8'h30;
    ff_ram[851] = 8'h10;
    ff_ram[852] = 8'h10;
    ff_ram[853] = 8'h10;
    ff_ram[854] = 8'h90;
    ff_ram[855] = 8'h60;
    ff_ram[856] = 8'h40;
    ff_ram[857] = 8'h40;
    ff_ram[858] = 8'h48;
    ff_ram[859] = 8'h50;
    ff_ram[860] = 8'h60;
    ff_ram[861] = 8'h50;
    ff_ram[862] = 8'h48;
    ff_ram[863] = 8'h00;
    ff_ram[864] = 8'h60;
    ff_ram[865] = 8'h20;
    ff_ram[866] = 8'h20;
    ff_ram[867] = 8'h20;
    ff_ram[868] = 8'h20;
    ff_ram[869] = 8'h20;
    ff_ram[870] = 8'h70;
    ff_ram[871] = 8'h00;
    ff_ram[872] = 8'h00;
    ff_ram[873] = 8'h00;
    ff_ram[874] = 8'hD0;
    ff_ram[875] = 8'hA8;
    ff_ram[876] = 8'hA8;
    ff_ram[877] = 8'hA8;
    ff_ram[878] = 8'hA8;
    ff_ram[879] = 8'h00;
    ff_ram[880] = 8'h00;
    ff_ram[881] = 8'h00;
    ff_ram[882] = 8'hB0;
    ff_ram[883] = 8'hC8;
    ff_ram[884] = 8'h88;
    ff_ram[885] = 8'h88;
    ff_ram[886] = 8'h88;
    ff_ram[887] = 8'h00;
    ff_ram[888] = 8'h00;
    ff_ram[889] = 8'h00;
    ff_ram[890] = 8'h70;
    ff_ram[891] = 8'h88;
    ff_ram[892] = 8'h88;
    ff_ram[893] = 8'h88;
    ff_ram[894] = 8'h70;
    ff_ram[895] = 8'h00;
    ff_ram[896] = 8'h00;
    ff_ram[897] = 8'h00;
    ff_ram[898] = 8'hB0;
    ff_ram[899] = 8'hC8;
    ff_ram[900] = 8'hC8;
    ff_ram[901] = 8'hB0;
    ff_ram[902] = 8'h80;
    ff_ram[903] = 8'h80;
    ff_ram[904] = 8'h00;
    ff_ram[905] = 8'h00;
    ff_ram[906] = 8'h68;
    ff_ram[907] = 8'h98;
    ff_ram[908] = 8'h98;
    ff_ram[909] = 8'h68;
    ff_ram[910] = 8'h08;
    ff_ram[911] = 8'h08;
    ff_ram[912] = 8'h00;
    ff_ram[913] = 8'h00;
    ff_ram[914] = 8'hB0;
    ff_ram[915] = 8'hC8;
    ff_ram[916] = 8'h80;
    ff_ram[917] = 8'h80;
    ff_ram[918] = 8'h80;
    ff_ram[919] = 8'h00;
    ff_ram[920] = 8'h00;
    ff_ram[921] = 8'h00;
    ff_ram[922] = 8'h78;
    ff_ram[923] = 8'h80;
    ff_ram[924] = 8'hF0;
    ff_ram[925] = 8'h08;
    ff_ram[926] = 8'hF0;
    ff_ram[927] = 8'h00;
    ff_ram[928] = 8'h40;
    ff_ram[929] = 8'h40;
    ff_ram[930] = 8'hF0;
    ff_ram[931] = 8'h40;
    ff_ram[932] = 8'h40;
    ff_ram[933] = 8'h48;
    ff_ram[934] = 8'h30;
    ff_ram[935] = 8'h00;
    ff_ram[936] = 8'h00;
    ff_ram[937] = 8'h00;
    ff_ram[938] = 8'h90;
    ff_ram[939] = 8'h90;
    ff_ram[940] = 8'h90;
    ff_ram[941] = 8'h90;
    ff_ram[942] = 8'h68;
    ff_ram[943] = 8'h00;
    ff_ram[944] = 8'h00;
    ff_ram[945] = 8'h00;
    ff_ram[946] = 8'h88;
    ff_ram[947] = 8'h88;
    ff_ram[948] = 8'h88;
    ff_ram[949] = 8'h50;
    ff_ram[950] = 8'h20;
    ff_ram[951] = 8'h00;
    ff_ram[952] = 8'h00;
    ff_ram[953] = 8'h00;
    ff_ram[954] = 8'h88;
    ff_ram[955] = 8'hA8;
    ff_ram[956] = 8'hA8;
    ff_ram[957] = 8'hA8;
    ff_ram[958] = 8'h50;
    ff_ram[959] = 8'h00;
    ff_ram[960] = 8'h00;
    ff_ram[961] = 8'h00;
    ff_ram[962] = 8'h88;
    ff_ram[963] = 8'h50;
    ff_ram[964] = 8'h20;
    ff_ram[965] = 8'h50;
    ff_ram[966] = 8'h88;
    ff_ram[967] = 8'h00;
    ff_ram[968] = 8'h00;
    ff_ram[969] = 8'h00;
    ff_ram[970] = 8'h88;
    ff_ram[971] = 8'h88;
    ff_ram[972] = 8'h98;
    ff_ram[973] = 8'h68;
    ff_ram[974] = 8'h08;
    ff_ram[975] = 8'h70;
    ff_ram[976] = 8'h00;
    ff_ram[977] = 8'h00;
    ff_ram[978] = 8'hF8;
    ff_ram[979] = 8'h10;
    ff_ram[980] = 8'h20;
    ff_ram[981] = 8'h40;
    ff_ram[982] = 8'hF8;
    ff_ram[983] = 8'h00;
    ff_ram[984] = 8'h18;
    ff_ram[985] = 8'h20;
    ff_ram[986] = 8'h20;
    ff_ram[987] = 8'h40;
    ff_ram[988] = 8'h20;
    ff_ram[989] = 8'h20;
    ff_ram[990] = 8'h18;
    ff_ram[991] = 8'h00;
    ff_ram[992] = 8'h20;
    ff_ram[993] = 8'h20;
    ff_ram[994] = 8'h20;
    ff_ram[995] = 8'h00;
    ff_ram[996] = 8'h20;
    ff_ram[997] = 8'h20;
    ff_ram[998] = 8'h20;
    ff_ram[999] = 8'h00;
    ff_ram[1000] = 8'hC0;
    ff_ram[1001] = 8'h20;
    ff_ram[1002] = 8'h20;
    ff_ram[1003] = 8'h10;
    ff_ram[1004] = 8'h20;
    ff_ram[1005] = 8'h20;
    ff_ram[1006] = 8'hC0;
    ff_ram[1007] = 8'h00;
    ff_ram[1008] = 8'h40;
    ff_ram[1009] = 8'hA8;
    ff_ram[1010] = 8'h10;
    ff_ram[1011] = 8'h00;
    ff_ram[1012] = 8'h00;
    ff_ram[1013] = 8'h00;
    ff_ram[1014] = 8'h00;
    ff_ram[1015] = 8'h00;
    ff_ram[1016] = 8'h00;
    ff_ram[1017] = 8'h00;
    ff_ram[1018] = 8'h00;
    ff_ram[1019] = 8'h00;
    ff_ram[1020] = 8'h00;
    ff_ram[1021] = 8'h00;
    ff_ram[1022] = 8'h00;
    ff_ram[1023] = 8'h00;
    ff_ram[1024] = 8'h10;
    ff_ram[1025] = 8'h38;
    ff_ram[1026] = 8'h7C;
    ff_ram[1027] = 8'hFE;
    ff_ram[1028] = 8'hFE;
    ff_ram[1029] = 8'h38;
    ff_ram[1030] = 8'h7C;
    ff_ram[1031] = 8'h00;
    ff_ram[1032] = 8'h6C;
    ff_ram[1033] = 8'hFE;
    ff_ram[1034] = 8'hFE;
    ff_ram[1035] = 8'hFE;
    ff_ram[1036] = 8'h7C;
    ff_ram[1037] = 8'h38;
    ff_ram[1038] = 8'h10;
    ff_ram[1039] = 8'h00;
    ff_ram[1040] = 8'h38;
    ff_ram[1041] = 8'h38;
    ff_ram[1042] = 8'hFE;
    ff_ram[1043] = 8'hFE;
    ff_ram[1044] = 8'hD6;
    ff_ram[1045] = 8'h10;
    ff_ram[1046] = 8'h7C;
    ff_ram[1047] = 8'h00;
    ff_ram[1048] = 8'h10;
    ff_ram[1049] = 8'h38;
    ff_ram[1050] = 8'h7C;
    ff_ram[1051] = 8'hFE;
    ff_ram[1052] = 8'h7C;
    ff_ram[1053] = 8'h38;
    ff_ram[1054] = 8'h10;
    ff_ram[1055] = 8'h00;
    ff_ram[1056] = 8'h00;
    ff_ram[1057] = 8'h78;
    ff_ram[1058] = 8'h84;
    ff_ram[1059] = 8'h84;
    ff_ram[1060] = 8'h84;
    ff_ram[1061] = 8'h84;
    ff_ram[1062] = 8'h78;
    ff_ram[1063] = 8'h00;
    ff_ram[1064] = 8'h00;
    ff_ram[1065] = 8'h78;
    ff_ram[1066] = 8'hFC;
    ff_ram[1067] = 8'hFC;
    ff_ram[1068] = 8'hFC;
    ff_ram[1069] = 8'hFC;
    ff_ram[1070] = 8'h78;
    ff_ram[1071] = 8'h00;
    ff_ram[1072] = 8'h20;
    ff_ram[1073] = 8'hF0;
    ff_ram[1074] = 8'h4C;
    ff_ram[1075] = 8'h70;
    ff_ram[1076] = 8'hA8;
    ff_ram[1077] = 8'h40;
    ff_ram[1078] = 8'h3C;
    ff_ram[1079] = 8'h00;
    ff_ram[1080] = 8'h00;
    ff_ram[1081] = 8'h20;
    ff_ram[1082] = 8'h78;
    ff_ram[1083] = 8'h20;
    ff_ram[1084] = 8'h78;
    ff_ram[1085] = 8'hB4;
    ff_ram[1086] = 8'h64;
    ff_ram[1087] = 8'h00;
    ff_ram[1088] = 8'h00;
    ff_ram[1089] = 8'h00;
    ff_ram[1090] = 8'h88;
    ff_ram[1091] = 8'h84;
    ff_ram[1092] = 8'h84;
    ff_ram[1093] = 8'h84;
    ff_ram[1094] = 8'h40;
    ff_ram[1095] = 8'h00;
    ff_ram[1096] = 8'h00;
    ff_ram[1097] = 8'h70;
    ff_ram[1098] = 8'h00;
    ff_ram[1099] = 8'h70;
    ff_ram[1100] = 8'h88;
    ff_ram[1101] = 8'h08;
    ff_ram[1102] = 8'h30;
    ff_ram[1103] = 8'h00;
    ff_ram[1104] = 8'h00;
    ff_ram[1105] = 8'h70;
    ff_ram[1106] = 8'h00;
    ff_ram[1107] = 8'hF0;
    ff_ram[1108] = 8'h20;
    ff_ram[1109] = 8'h60;
    ff_ram[1110] = 8'h98;
    ff_ram[1111] = 8'h00;
    ff_ram[1112] = 8'h00;
    ff_ram[1113] = 8'h20;
    ff_ram[1114] = 8'hF8;
    ff_ram[1115] = 8'h24;
    ff_ram[1116] = 8'h78;
    ff_ram[1117] = 8'hA4;
    ff_ram[1118] = 8'h68;
    ff_ram[1119] = 8'h00;
    ff_ram[1120] = 8'h00;
    ff_ram[1121] = 8'h90;
    ff_ram[1122] = 8'h58;
    ff_ram[1123] = 8'h64;
    ff_ram[1124] = 8'hA8;
    ff_ram[1125] = 8'h20;
    ff_ram[1126] = 8'h10;
    ff_ram[1127] = 8'h00;
    ff_ram[1128] = 8'h00;
    ff_ram[1129] = 8'h10;
    ff_ram[1130] = 8'hB8;
    ff_ram[1131] = 8'hD4;
    ff_ram[1132] = 8'h94;
    ff_ram[1133] = 8'h18;
    ff_ram[1134] = 8'h20;
    ff_ram[1135] = 8'h00;
    ff_ram[1136] = 8'h00;
    ff_ram[1137] = 8'h10;
    ff_ram[1138] = 8'h1C;
    ff_ram[1139] = 8'h10;
    ff_ram[1140] = 8'h70;
    ff_ram[1141] = 8'h98;
    ff_ram[1142] = 8'h74;
    ff_ram[1143] = 8'h00;
    ff_ram[1144] = 8'h00;
    ff_ram[1145] = 8'h00;
    ff_ram[1146] = 8'h00;
    ff_ram[1147] = 8'h78;
    ff_ram[1148] = 8'h04;
    ff_ram[1149] = 8'h04;
    ff_ram[1150] = 8'h38;
    ff_ram[1151] = 8'h00;
    ff_ram[1152] = 8'h00;
    ff_ram[1153] = 8'h00;
    ff_ram[1154] = 8'h00;
    ff_ram[1155] = 8'h00;
    ff_ram[1156] = 8'h00;
    ff_ram[1157] = 8'h00;
    ff_ram[1158] = 8'h00;
    ff_ram[1159] = 8'h00;
    ff_ram[1160] = 8'h20;
    ff_ram[1161] = 8'h7C;
    ff_ram[1162] = 8'h20;
    ff_ram[1163] = 8'h7C;
    ff_ram[1164] = 8'hAA;
    ff_ram[1165] = 8'h92;
    ff_ram[1166] = 8'h64;
    ff_ram[1167] = 8'h00;
    ff_ram[1168] = 8'h00;
    ff_ram[1169] = 8'h84;
    ff_ram[1170] = 8'h82;
    ff_ram[1171] = 8'h82;
    ff_ram[1172] = 8'h82;
    ff_ram[1173] = 8'h80;
    ff_ram[1174] = 8'h40;
    ff_ram[1175] = 8'h00;
    ff_ram[1176] = 8'h38;
    ff_ram[1177] = 8'h00;
    ff_ram[1178] = 8'h38;
    ff_ram[1179] = 8'h44;
    ff_ram[1180] = 8'h04;
    ff_ram[1181] = 8'h08;
    ff_ram[1182] = 8'h30;
    ff_ram[1183] = 8'h00;
    ff_ram[1184] = 8'h70;
    ff_ram[1185] = 8'h00;
    ff_ram[1186] = 8'hF8;
    ff_ram[1187] = 8'h10;
    ff_ram[1188] = 8'h20;
    ff_ram[1189] = 8'h60;
    ff_ram[1190] = 8'h9C;
    ff_ram[1191] = 8'h00;
    ff_ram[1192] = 8'h24;
    ff_ram[1193] = 8'hFA;
    ff_ram[1194] = 8'h20;
    ff_ram[1195] = 8'h7C;
    ff_ram[1196] = 8'hA2;
    ff_ram[1197] = 8'hA2;
    ff_ram[1198] = 8'h44;
    ff_ram[1199] = 8'h00;
    ff_ram[1200] = 8'h40;
    ff_ram[1201] = 8'h44;
    ff_ram[1202] = 8'hF2;
    ff_ram[1203] = 8'h4A;
    ff_ram[1204] = 8'h48;
    ff_ram[1205] = 8'h88;
    ff_ram[1206] = 8'h30;
    ff_ram[1207] = 8'h00;
    ff_ram[1208] = 8'h20;
    ff_ram[1209] = 8'hFC;
    ff_ram[1210] = 8'h10;
    ff_ram[1211] = 8'hFC;
    ff_ram[1212] = 8'h08;
    ff_ram[1213] = 8'h80;
    ff_ram[1214] = 8'h78;
    ff_ram[1215] = 8'h00;
    ff_ram[1216] = 8'h08;
    ff_ram[1217] = 8'h10;
    ff_ram[1218] = 8'h20;
    ff_ram[1219] = 8'h40;
    ff_ram[1220] = 8'h20;
    ff_ram[1221] = 8'h10;
    ff_ram[1222] = 8'h08;
    ff_ram[1223] = 8'h00;
    ff_ram[1224] = 8'h04;
    ff_ram[1225] = 8'h84;
    ff_ram[1226] = 8'h9E;
    ff_ram[1227] = 8'h84;
    ff_ram[1228] = 8'h84;
    ff_ram[1229] = 8'h84;
    ff_ram[1230] = 8'h48;
    ff_ram[1231] = 8'h00;
    ff_ram[1232] = 8'h78;
    ff_ram[1233] = 8'h04;
    ff_ram[1234] = 8'h00;
    ff_ram[1235] = 8'h00;
    ff_ram[1236] = 8'h00;
    ff_ram[1237] = 8'h80;
    ff_ram[1238] = 8'h7C;
    ff_ram[1239] = 8'h00;
    ff_ram[1240] = 8'h10;
    ff_ram[1241] = 8'hFE;
    ff_ram[1242] = 8'h08;
    ff_ram[1243] = 8'h04;
    ff_ram[1244] = 8'h04;
    ff_ram[1245] = 8'h80;
    ff_ram[1246] = 8'h78;
    ff_ram[1247] = 8'h00;
    ff_ram[1248] = 8'h80;
    ff_ram[1249] = 8'h80;
    ff_ram[1250] = 8'h80;
    ff_ram[1251] = 8'h80;
    ff_ram[1252] = 8'h84;
    ff_ram[1253] = 8'h88;
    ff_ram[1254] = 8'h70;
    ff_ram[1255] = 8'h00;
    ff_ram[1256] = 8'h08;
    ff_ram[1257] = 8'hFE;
    ff_ram[1258] = 8'h38;
    ff_ram[1259] = 8'h48;
    ff_ram[1260] = 8'h38;
    ff_ram[1261] = 8'h08;
    ff_ram[1262] = 8'h10;
    ff_ram[1263] = 8'h00;
    ff_ram[1264] = 8'h44;
    ff_ram[1265] = 8'h44;
    ff_ram[1266] = 8'hFE;
    ff_ram[1267] = 8'h44;
    ff_ram[1268] = 8'h48;
    ff_ram[1269] = 8'h40;
    ff_ram[1270] = 8'h3C;
    ff_ram[1271] = 8'h00;
    ff_ram[1272] = 8'h44;
    ff_ram[1273] = 8'h28;
    ff_ram[1274] = 8'hFE;
    ff_ram[1275] = 8'h20;
    ff_ram[1276] = 8'h40;
    ff_ram[1277] = 8'h40;
    ff_ram[1278] = 8'h3C;
    ff_ram[1279] = 8'h00;
    ff_ram[1280] = 8'h00;
    ff_ram[1281] = 8'h00;
    ff_ram[1282] = 8'h00;
    ff_ram[1283] = 8'h00;
    ff_ram[1284] = 8'h00;
    ff_ram[1285] = 8'h00;
    ff_ram[1286] = 8'h00;
    ff_ram[1287] = 8'h00;
    ff_ram[1288] = 8'h00;
    ff_ram[1289] = 8'h00;
    ff_ram[1290] = 8'h00;
    ff_ram[1291] = 8'h00;
    ff_ram[1292] = 8'h60;
    ff_ram[1293] = 8'h90;
    ff_ram[1294] = 8'h60;
    ff_ram[1295] = 8'h00;
    ff_ram[1296] = 8'h38;
    ff_ram[1297] = 8'h20;
    ff_ram[1298] = 8'h20;
    ff_ram[1299] = 8'h20;
    ff_ram[1300] = 8'h00;
    ff_ram[1301] = 8'h00;
    ff_ram[1302] = 8'h00;
    ff_ram[1303] = 8'h00;
    ff_ram[1304] = 8'h00;
    ff_ram[1305] = 8'h00;
    ff_ram[1306] = 8'h00;
    ff_ram[1307] = 8'h20;
    ff_ram[1308] = 8'h20;
    ff_ram[1309] = 8'h20;
    ff_ram[1310] = 8'hE0;
    ff_ram[1311] = 8'h00;
    ff_ram[1312] = 8'h00;
    ff_ram[1313] = 8'h00;
    ff_ram[1314] = 8'h00;
    ff_ram[1315] = 8'h00;
    ff_ram[1316] = 8'h80;
    ff_ram[1317] = 8'h40;
    ff_ram[1318] = 8'h20;
    ff_ram[1319] = 8'h00;
    ff_ram[1320] = 8'h00;
    ff_ram[1321] = 8'h00;
    ff_ram[1322] = 8'h00;
    ff_ram[1323] = 8'h30;
    ff_ram[1324] = 8'h30;
    ff_ram[1325] = 8'h00;
    ff_ram[1326] = 8'h00;
    ff_ram[1327] = 8'h00;
    ff_ram[1328] = 8'hF8;
    ff_ram[1329] = 8'h08;
    ff_ram[1330] = 8'hF8;
    ff_ram[1331] = 8'h08;
    ff_ram[1332] = 8'h10;
    ff_ram[1333] = 8'h20;
    ff_ram[1334] = 8'h40;
    ff_ram[1335] = 8'h00;
    ff_ram[1336] = 8'h00;
    ff_ram[1337] = 8'h00;
    ff_ram[1338] = 8'hF0;
    ff_ram[1339] = 8'h10;
    ff_ram[1340] = 8'h60;
    ff_ram[1341] = 8'h40;
    ff_ram[1342] = 8'h80;
    ff_ram[1343] = 8'h00;
    ff_ram[1344] = 8'h00;
    ff_ram[1345] = 8'h10;
    ff_ram[1346] = 8'h20;
    ff_ram[1347] = 8'h60;
    ff_ram[1348] = 8'hA0;
    ff_ram[1349] = 8'h20;
    ff_ram[1350] = 8'h20;
    ff_ram[1351] = 8'h00;
    ff_ram[1352] = 8'h00;
    ff_ram[1353] = 8'h20;
    ff_ram[1354] = 8'hF0;
    ff_ram[1355] = 8'h90;
    ff_ram[1356] = 8'h10;
    ff_ram[1357] = 8'h20;
    ff_ram[1358] = 8'h40;
    ff_ram[1359] = 8'h00;
    ff_ram[1360] = 8'h00;
    ff_ram[1361] = 8'h00;
    ff_ram[1362] = 8'hF0;
    ff_ram[1363] = 8'h20;
    ff_ram[1364] = 8'h20;
    ff_ram[1365] = 8'h20;
    ff_ram[1366] = 8'hF0;
    ff_ram[1367] = 8'h00;
    ff_ram[1368] = 8'h00;
    ff_ram[1369] = 8'h20;
    ff_ram[1370] = 8'hF0;
    ff_ram[1371] = 8'h60;
    ff_ram[1372] = 8'hA0;
    ff_ram[1373] = 8'hA0;
    ff_ram[1374] = 8'h20;
    ff_ram[1375] = 8'h00;
    ff_ram[1376] = 8'h00;
    ff_ram[1377] = 8'h40;
    ff_ram[1378] = 8'hF8;
    ff_ram[1379] = 8'h48;
    ff_ram[1380] = 8'h50;
    ff_ram[1381] = 8'h40;
    ff_ram[1382] = 8'h40;
    ff_ram[1383] = 8'h00;
    ff_ram[1384] = 8'h00;
    ff_ram[1385] = 8'h00;
    ff_ram[1386] = 8'h70;
    ff_ram[1387] = 8'h10;
    ff_ram[1388] = 8'h10;
    ff_ram[1389] = 8'h10;
    ff_ram[1390] = 8'hF8;
    ff_ram[1391] = 8'h00;
    ff_ram[1392] = 8'h00;
    ff_ram[1393] = 8'h00;
    ff_ram[1394] = 8'hF0;
    ff_ram[1395] = 8'h10;
    ff_ram[1396] = 8'hF0;
    ff_ram[1397] = 8'h10;
    ff_ram[1398] = 8'hF0;
    ff_ram[1399] = 8'h00;
    ff_ram[1400] = 8'h00;
    ff_ram[1401] = 8'h00;
    ff_ram[1402] = 8'hA8;
    ff_ram[1403] = 8'hA8;
    ff_ram[1404] = 8'h08;
    ff_ram[1405] = 8'h10;
    ff_ram[1406] = 8'h20;
    ff_ram[1407] = 8'h00;
    ff_ram[1408] = 8'h00;
    ff_ram[1409] = 8'h00;
    ff_ram[1410] = 8'h80;
    ff_ram[1411] = 8'h7C;
    ff_ram[1412] = 8'h00;
    ff_ram[1413] = 8'h00;
    ff_ram[1414] = 8'h00;
    ff_ram[1415] = 8'h00;
    ff_ram[1416] = 8'hF8;
    ff_ram[1417] = 8'h08;
    ff_ram[1418] = 8'h28;
    ff_ram[1419] = 8'h30;
    ff_ram[1420] = 8'h20;
    ff_ram[1421] = 8'h20;
    ff_ram[1422] = 8'h40;
    ff_ram[1423] = 8'h00;
    ff_ram[1424] = 8'h08;
    ff_ram[1425] = 8'h10;
    ff_ram[1426] = 8'h20;
    ff_ram[1427] = 8'h60;
    ff_ram[1428] = 8'hA0;
    ff_ram[1429] = 8'h20;
    ff_ram[1430] = 8'h20;
    ff_ram[1431] = 8'h00;
    ff_ram[1432] = 8'h20;
    ff_ram[1433] = 8'hF8;
    ff_ram[1434] = 8'h88;
    ff_ram[1435] = 8'h88;
    ff_ram[1436] = 8'h08;
    ff_ram[1437] = 8'h10;
    ff_ram[1438] = 8'h20;
    ff_ram[1439] = 8'h00;
    ff_ram[1440] = 8'h00;
    ff_ram[1441] = 8'hF8;
    ff_ram[1442] = 8'h20;
    ff_ram[1443] = 8'h20;
    ff_ram[1444] = 8'h20;
    ff_ram[1445] = 8'h20;
    ff_ram[1446] = 8'hF8;
    ff_ram[1447] = 8'h00;
    ff_ram[1448] = 8'h10;
    ff_ram[1449] = 8'hF8;
    ff_ram[1450] = 8'h10;
    ff_ram[1451] = 8'h30;
    ff_ram[1452] = 8'h50;
    ff_ram[1453] = 8'h90;
    ff_ram[1454] = 8'h10;
    ff_ram[1455] = 8'h00;
    ff_ram[1456] = 8'h20;
    ff_ram[1457] = 8'hF8;
    ff_ram[1458] = 8'h28;
    ff_ram[1459] = 8'h28;
    ff_ram[1460] = 8'h28;
    ff_ram[1461] = 8'h48;
    ff_ram[1462] = 8'h88;
    ff_ram[1463] = 8'h00;
    ff_ram[1464] = 8'h20;
    ff_ram[1465] = 8'hF8;
    ff_ram[1466] = 8'h20;
    ff_ram[1467] = 8'hF8;
    ff_ram[1468] = 8'h20;
    ff_ram[1469] = 8'h20;
    ff_ram[1470] = 8'h20;
    ff_ram[1471] = 8'h00;
    ff_ram[1472] = 8'h78;
    ff_ram[1473] = 8'h48;
    ff_ram[1474] = 8'h88;
    ff_ram[1475] = 8'h08;
    ff_ram[1476] = 8'h08;
    ff_ram[1477] = 8'h10;
    ff_ram[1478] = 8'h20;
    ff_ram[1479] = 8'h00;
    ff_ram[1480] = 8'h40;
    ff_ram[1481] = 8'h78;
    ff_ram[1482] = 8'h50;
    ff_ram[1483] = 8'h90;
    ff_ram[1484] = 8'h10;
    ff_ram[1485] = 8'h10;
    ff_ram[1486] = 8'h20;
    ff_ram[1487] = 8'h00;
    ff_ram[1488] = 8'h00;
    ff_ram[1489] = 8'hF8;
    ff_ram[1490] = 8'h08;
    ff_ram[1491] = 8'h08;
    ff_ram[1492] = 8'h08;
    ff_ram[1493] = 8'h08;
    ff_ram[1494] = 8'hF8;
    ff_ram[1495] = 8'h00;
    ff_ram[1496] = 8'h50;
    ff_ram[1497] = 8'hF8;
    ff_ram[1498] = 8'h50;
    ff_ram[1499] = 8'h50;
    ff_ram[1500] = 8'h10;
    ff_ram[1501] = 8'h10;
    ff_ram[1502] = 8'h20;
    ff_ram[1503] = 8'h00;
    ff_ram[1504] = 8'h00;
    ff_ram[1505] = 8'hC0;
    ff_ram[1506] = 8'h08;
    ff_ram[1507] = 8'hC8;
    ff_ram[1508] = 8'h08;
    ff_ram[1509] = 8'h10;
    ff_ram[1510] = 8'hE0;
    ff_ram[1511] = 8'h00;
    ff_ram[1512] = 8'h00;
    ff_ram[1513] = 8'hF8;
    ff_ram[1514] = 8'h08;
    ff_ram[1515] = 8'h10;
    ff_ram[1516] = 8'h20;
    ff_ram[1517] = 8'h50;
    ff_ram[1518] = 8'h88;
    ff_ram[1519] = 8'h00;
    ff_ram[1520] = 8'h40;
    ff_ram[1521] = 8'hF8;
    ff_ram[1522] = 8'h48;
    ff_ram[1523] = 8'h50;
    ff_ram[1524] = 8'h40;
    ff_ram[1525] = 8'h40;
    ff_ram[1526] = 8'h38;
    ff_ram[1527] = 8'h00;
    ff_ram[1528] = 8'h88;
    ff_ram[1529] = 8'h88;
    ff_ram[1530] = 8'h48;
    ff_ram[1531] = 8'h08;
    ff_ram[1532] = 8'h10;
    ff_ram[1533] = 8'h20;
    ff_ram[1534] = 8'h40;
    ff_ram[1535] = 8'h00;
    ff_ram[1536] = 8'h78;
    ff_ram[1537] = 8'h48;
    ff_ram[1538] = 8'h78;
    ff_ram[1539] = 8'h88;
    ff_ram[1540] = 8'h08;
    ff_ram[1541] = 8'h10;
    ff_ram[1542] = 8'h20;
    ff_ram[1543] = 8'h00;
    ff_ram[1544] = 8'h10;
    ff_ram[1545] = 8'hE0;
    ff_ram[1546] = 8'h20;
    ff_ram[1547] = 8'hF8;
    ff_ram[1548] = 8'h20;
    ff_ram[1549] = 8'h20;
    ff_ram[1550] = 8'h40;
    ff_ram[1551] = 8'h00;
    ff_ram[1552] = 8'hA8;
    ff_ram[1553] = 8'hA8;
    ff_ram[1554] = 8'hA8;
    ff_ram[1555] = 8'h08;
    ff_ram[1556] = 8'h08;
    ff_ram[1557] = 8'h10;
    ff_ram[1558] = 8'h20;
    ff_ram[1559] = 8'h00;
    ff_ram[1560] = 8'h70;
    ff_ram[1561] = 8'h00;
    ff_ram[1562] = 8'hF8;
    ff_ram[1563] = 8'h20;
    ff_ram[1564] = 8'h20;
    ff_ram[1565] = 8'h20;
    ff_ram[1566] = 8'h40;
    ff_ram[1567] = 8'h00;
    ff_ram[1568] = 8'h40;
    ff_ram[1569] = 8'h40;
    ff_ram[1570] = 8'h60;
    ff_ram[1571] = 8'h50;
    ff_ram[1572] = 8'h48;
    ff_ram[1573] = 8'h40;
    ff_ram[1574] = 8'h40;
    ff_ram[1575] = 8'h00;
    ff_ram[1576] = 8'h20;
    ff_ram[1577] = 8'hF8;
    ff_ram[1578] = 8'h20;
    ff_ram[1579] = 8'h20;
    ff_ram[1580] = 8'h20;
    ff_ram[1581] = 8'h20;
    ff_ram[1582] = 8'h40;
    ff_ram[1583] = 8'h00;
    ff_ram[1584] = 8'h00;
    ff_ram[1585] = 8'h70;
    ff_ram[1586] = 8'h00;
    ff_ram[1587] = 8'h00;
    ff_ram[1588] = 8'h00;
    ff_ram[1589] = 8'h00;
    ff_ram[1590] = 8'hF8;
    ff_ram[1591] = 8'h00;
    ff_ram[1592] = 8'h00;
    ff_ram[1593] = 8'hF8;
    ff_ram[1594] = 8'h08;
    ff_ram[1595] = 8'hD0;
    ff_ram[1596] = 8'h20;
    ff_ram[1597] = 8'h50;
    ff_ram[1598] = 8'h88;
    ff_ram[1599] = 8'h00;
    ff_ram[1600] = 8'h20;
    ff_ram[1601] = 8'hF8;
    ff_ram[1602] = 8'h08;
    ff_ram[1603] = 8'h30;
    ff_ram[1604] = 8'hE8;
    ff_ram[1605] = 8'h20;
    ff_ram[1606] = 8'h20;
    ff_ram[1607] = 8'h00;
    ff_ram[1608] = 8'h08;
    ff_ram[1609] = 8'h08;
    ff_ram[1610] = 8'h08;
    ff_ram[1611] = 8'h10;
    ff_ram[1612] = 8'h20;
    ff_ram[1613] = 8'h40;
    ff_ram[1614] = 8'h80;
    ff_ram[1615] = 8'h00;
    ff_ram[1616] = 8'h20;
    ff_ram[1617] = 8'h10;
    ff_ram[1618] = 8'h48;
    ff_ram[1619] = 8'h48;
    ff_ram[1620] = 8'h48;
    ff_ram[1621] = 8'h48;
    ff_ram[1622] = 8'h88;
    ff_ram[1623] = 8'h00;
    ff_ram[1624] = 8'h80;
    ff_ram[1625] = 8'h80;
    ff_ram[1626] = 8'hF8;
    ff_ram[1627] = 8'h80;
    ff_ram[1628] = 8'h80;
    ff_ram[1629] = 8'h80;
    ff_ram[1630] = 8'h78;
    ff_ram[1631] = 8'h00;
    ff_ram[1632] = 8'hF8;
    ff_ram[1633] = 8'h08;
    ff_ram[1634] = 8'h08;
    ff_ram[1635] = 8'h08;
    ff_ram[1636] = 8'h10;
    ff_ram[1637] = 8'h20;
    ff_ram[1638] = 8'h40;
    ff_ram[1639] = 8'h00;
    ff_ram[1640] = 8'h00;
    ff_ram[1641] = 8'h40;
    ff_ram[1642] = 8'hA0;
    ff_ram[1643] = 8'h10;
    ff_ram[1644] = 8'h08;
    ff_ram[1645] = 8'h08;
    ff_ram[1646] = 8'h00;
    ff_ram[1647] = 8'h00;
    ff_ram[1648] = 8'h20;
    ff_ram[1649] = 8'hF8;
    ff_ram[1650] = 8'h20;
    ff_ram[1651] = 8'h20;
    ff_ram[1652] = 8'hA8;
    ff_ram[1653] = 8'hA8;
    ff_ram[1654] = 8'h20;
    ff_ram[1655] = 8'h00;
    ff_ram[1656] = 8'h00;
    ff_ram[1657] = 8'hF8;
    ff_ram[1658] = 8'h08;
    ff_ram[1659] = 8'h08;
    ff_ram[1660] = 8'h50;
    ff_ram[1661] = 8'h20;
    ff_ram[1662] = 8'h10;
    ff_ram[1663] = 8'h00;
    ff_ram[1664] = 8'hF0;
    ff_ram[1665] = 8'h00;
    ff_ram[1666] = 8'h60;
    ff_ram[1667] = 8'h00;
    ff_ram[1668] = 8'h00;
    ff_ram[1669] = 8'hF0;
    ff_ram[1670] = 8'h08;
    ff_ram[1671] = 8'h00;
    ff_ram[1672] = 8'h10;
    ff_ram[1673] = 8'h20;
    ff_ram[1674] = 8'h40;
    ff_ram[1675] = 8'h80;
    ff_ram[1676] = 8'h90;
    ff_ram[1677] = 8'h88;
    ff_ram[1678] = 8'hF8;
    ff_ram[1679] = 8'h00;
    ff_ram[1680] = 8'h08;
    ff_ram[1681] = 8'h08;
    ff_ram[1682] = 8'h08;
    ff_ram[1683] = 8'h50;
    ff_ram[1684] = 8'h20;
    ff_ram[1685] = 8'h50;
    ff_ram[1686] = 8'h80;
    ff_ram[1687] = 8'h00;
    ff_ram[1688] = 8'h78;
    ff_ram[1689] = 8'h20;
    ff_ram[1690] = 8'hF8;
    ff_ram[1691] = 8'h20;
    ff_ram[1692] = 8'h20;
    ff_ram[1693] = 8'h20;
    ff_ram[1694] = 8'h18;
    ff_ram[1695] = 8'h00;
    ff_ram[1696] = 8'h40;
    ff_ram[1697] = 8'hF8;
    ff_ram[1698] = 8'h48;
    ff_ram[1699] = 8'h48;
    ff_ram[1700] = 8'h50;
    ff_ram[1701] = 8'h40;
    ff_ram[1702] = 8'h40;
    ff_ram[1703] = 8'h00;
    ff_ram[1704] = 8'h00;
    ff_ram[1705] = 8'h70;
    ff_ram[1706] = 8'h10;
    ff_ram[1707] = 8'h10;
    ff_ram[1708] = 8'h10;
    ff_ram[1709] = 8'h10;
    ff_ram[1710] = 8'hF8;
    ff_ram[1711] = 8'h00;
    ff_ram[1712] = 8'h00;
    ff_ram[1713] = 8'hF8;
    ff_ram[1714] = 8'h08;
    ff_ram[1715] = 8'hF8;
    ff_ram[1716] = 8'h08;
    ff_ram[1717] = 8'h08;
    ff_ram[1718] = 8'hF8;
    ff_ram[1719] = 8'h00;
    ff_ram[1720] = 8'h70;
    ff_ram[1721] = 8'h00;
    ff_ram[1722] = 8'hF8;
    ff_ram[1723] = 8'h08;
    ff_ram[1724] = 8'h08;
    ff_ram[1725] = 8'h10;
    ff_ram[1726] = 8'h20;
    ff_ram[1727] = 8'h00;
    ff_ram[1728] = 8'h48;
    ff_ram[1729] = 8'h48;
    ff_ram[1730] = 8'h48;
    ff_ram[1731] = 8'h48;
    ff_ram[1732] = 8'h48;
    ff_ram[1733] = 8'h10;
    ff_ram[1734] = 8'h20;
    ff_ram[1735] = 8'h00;
    ff_ram[1736] = 8'h10;
    ff_ram[1737] = 8'h50;
    ff_ram[1738] = 8'h50;
    ff_ram[1739] = 8'h50;
    ff_ram[1740] = 8'h50;
    ff_ram[1741] = 8'h58;
    ff_ram[1742] = 8'h90;
    ff_ram[1743] = 8'h00;
    ff_ram[1744] = 8'h40;
    ff_ram[1745] = 8'h40;
    ff_ram[1746] = 8'h40;
    ff_ram[1747] = 8'h48;
    ff_ram[1748] = 8'h48;
    ff_ram[1749] = 8'h50;
    ff_ram[1750] = 8'h60;
    ff_ram[1751] = 8'h00;
    ff_ram[1752] = 8'h00;
    ff_ram[1753] = 8'hF8;
    ff_ram[1754] = 8'h88;
    ff_ram[1755] = 8'h88;
    ff_ram[1756] = 8'h88;
    ff_ram[1757] = 8'h88;
    ff_ram[1758] = 8'hF8;
    ff_ram[1759] = 8'h00;
    ff_ram[1760] = 8'hF8;
    ff_ram[1761] = 8'h88;
    ff_ram[1762] = 8'h88;
    ff_ram[1763] = 8'h08;
    ff_ram[1764] = 8'h08;
    ff_ram[1765] = 8'h10;
    ff_ram[1766] = 8'h20;
    ff_ram[1767] = 8'h00;
    ff_ram[1768] = 8'h00;
    ff_ram[1769] = 8'hC0;
    ff_ram[1770] = 8'h00;
    ff_ram[1771] = 8'h08;
    ff_ram[1772] = 8'h08;
    ff_ram[1773] = 8'h10;
    ff_ram[1774] = 8'hE0;
    ff_ram[1775] = 8'h00;
    ff_ram[1776] = 8'h90;
    ff_ram[1777] = 8'h48;
    ff_ram[1778] = 8'h00;
    ff_ram[1779] = 8'h00;
    ff_ram[1780] = 8'h00;
    ff_ram[1781] = 8'h00;
    ff_ram[1782] = 8'h00;
    ff_ram[1783] = 8'h00;
    ff_ram[1784] = 8'h60;
    ff_ram[1785] = 8'h90;
    ff_ram[1786] = 8'h60;
    ff_ram[1787] = 8'h00;
    ff_ram[1788] = 8'h00;
    ff_ram[1789] = 8'h00;
    ff_ram[1790] = 8'h00;
    ff_ram[1791] = 8'h00;
    ff_ram[1792] = 8'h20;
    ff_ram[1793] = 8'hF8;
    ff_ram[1794] = 8'h20;
    ff_ram[1795] = 8'h4E;
    ff_ram[1796] = 8'h40;
    ff_ram[1797] = 8'h90;
    ff_ram[1798] = 8'h8E;
    ff_ram[1799] = 8'h00;
    ff_ram[1800] = 8'h10;
    ff_ram[1801] = 8'hFE;
    ff_ram[1802] = 8'h20;
    ff_ram[1803] = 8'h78;
    ff_ram[1804] = 8'h04;
    ff_ram[1805] = 8'h04;
    ff_ram[1806] = 8'h78;
    ff_ram[1807] = 8'h00;
    ff_ram[1808] = 8'h00;
    ff_ram[1809] = 8'hFC;
    ff_ram[1810] = 8'h02;
    ff_ram[1811] = 8'h02;
    ff_ram[1812] = 8'h02;
    ff_ram[1813] = 8'h04;
    ff_ram[1814] = 8'h18;
    ff_ram[1815] = 8'h00;
    ff_ram[1816] = 8'hFE;
    ff_ram[1817] = 8'h08;
    ff_ram[1818] = 8'h10;
    ff_ram[1819] = 8'h20;
    ff_ram[1820] = 8'h20;
    ff_ram[1821] = 8'h20;
    ff_ram[1822] = 8'h1C;
    ff_ram[1823] = 8'h00;
    ff_ram[1824] = 8'h20;
    ff_ram[1825] = 8'h24;
    ff_ram[1826] = 8'h38;
    ff_ram[1827] = 8'h60;
    ff_ram[1828] = 8'h80;
    ff_ram[1829] = 8'h80;
    ff_ram[1830] = 8'h7C;
    ff_ram[1831] = 8'h00;
    ff_ram[1832] = 8'h2C;
    ff_ram[1833] = 8'hF2;
    ff_ram[1834] = 8'h44;
    ff_ram[1835] = 8'h44;
    ff_ram[1836] = 8'h9C;
    ff_ram[1837] = 8'h26;
    ff_ram[1838] = 8'h1C;
    ff_ram[1839] = 8'h00;
    ff_ram[1840] = 8'h00;
    ff_ram[1841] = 8'h9E;
    ff_ram[1842] = 8'h80;
    ff_ram[1843] = 8'h80;
    ff_ram[1844] = 8'h80;
    ff_ram[1845] = 8'h90;
    ff_ram[1846] = 8'h4E;
    ff_ram[1847] = 8'h00;
    ff_ram[1848] = 8'h48;
    ff_ram[1849] = 8'h48;
    ff_ram[1850] = 8'h7C;
    ff_ram[1851] = 8'hD2;
    ff_ram[1852] = 8'hB6;
    ff_ram[1853] = 8'hAA;
    ff_ram[1854] = 8'h4C;
    ff_ram[1855] = 8'h00;
    ff_ram[1856] = 8'h40;
    ff_ram[1857] = 8'h4C;
    ff_ram[1858] = 8'hD2;
    ff_ram[1859] = 8'h62;
    ff_ram[1860] = 8'h4E;
    ff_ram[1861] = 8'hD2;
    ff_ram[1862] = 8'h4E;
    ff_ram[1863] = 8'h00;
    ff_ram[1864] = 8'h00;
    ff_ram[1865] = 8'h38;
    ff_ram[1866] = 8'h54;
    ff_ram[1867] = 8'h92;
    ff_ram[1868] = 8'hA2;
    ff_ram[1869] = 8'hA2;
    ff_ram[1870] = 8'h44;
    ff_ram[1871] = 8'h00;
    ff_ram[1872] = 8'h04;
    ff_ram[1873] = 8'h9E;
    ff_ram[1874] = 8'h84;
    ff_ram[1875] = 8'h84;
    ff_ram[1876] = 8'h8C;
    ff_ram[1877] = 8'h96;
    ff_ram[1878] = 8'h4C;
    ff_ram[1879] = 8'h00;
    ff_ram[1880] = 8'h10;
    ff_ram[1881] = 8'hE4;
    ff_ram[1882] = 8'h26;
    ff_ram[1883] = 8'h44;
    ff_ram[1884] = 8'h44;
    ff_ram[1885] = 8'h48;
    ff_ram[1886] = 8'h30;
    ff_ram[1887] = 8'h00;
    ff_ram[1888] = 8'h20;
    ff_ram[1889] = 8'h10;
    ff_ram[1890] = 8'h00;
    ff_ram[1891] = 8'h20;
    ff_ram[1892] = 8'h14;
    ff_ram[1893] = 8'h52;
    ff_ram[1894] = 8'hB2;
    ff_ram[1895] = 8'h00;
    ff_ram[1896] = 8'h00;
    ff_ram[1897] = 8'h00;
    ff_ram[1898] = 8'h20;
    ff_ram[1899] = 8'h50;
    ff_ram[1900] = 8'h88;
    ff_ram[1901] = 8'h04;
    ff_ram[1902] = 8'h02;
    ff_ram[1903] = 8'h00;
    ff_ram[1904] = 8'h1E;
    ff_ram[1905] = 8'h84;
    ff_ram[1906] = 8'h9E;
    ff_ram[1907] = 8'h84;
    ff_ram[1908] = 8'h8C;
    ff_ram[1909] = 8'h96;
    ff_ram[1910] = 8'h4C;
    ff_ram[1911] = 8'h00;
    ff_ram[1912] = 8'h10;
    ff_ram[1913] = 8'hFC;
    ff_ram[1914] = 8'h10;
    ff_ram[1915] = 8'hFC;
    ff_ram[1916] = 8'h70;
    ff_ram[1917] = 8'h98;
    ff_ram[1918] = 8'h74;
    ff_ram[1919] = 8'h00;
    ff_ram[1920] = 8'h70;
    ff_ram[1921] = 8'h10;
    ff_ram[1922] = 8'h14;
    ff_ram[1923] = 8'h7E;
    ff_ram[1924] = 8'hA4;
    ff_ram[1925] = 8'hA4;
    ff_ram[1926] = 8'h48;
    ff_ram[1927] = 8'h00;
    ff_ram[1928] = 8'h20;
    ff_ram[1929] = 8'hF4;
    ff_ram[1930] = 8'h22;
    ff_ram[1931] = 8'h60;
    ff_ram[1932] = 8'hA2;
    ff_ram[1933] = 8'h62;
    ff_ram[1934] = 8'h1C;
    ff_ram[1935] = 8'h00;
    ff_ram[1936] = 8'h48;
    ff_ram[1937] = 8'h48;
    ff_ram[1938] = 8'h7C;
    ff_ram[1939] = 8'hAA;
    ff_ram[1940] = 8'h92;
    ff_ram[1941] = 8'hA2;
    ff_ram[1942] = 8'h44;
    ff_ram[1943] = 8'h00;
    ff_ram[1944] = 8'h20;
    ff_ram[1945] = 8'hF8;
    ff_ram[1946] = 8'h20;
    ff_ram[1947] = 8'hF8;
    ff_ram[1948] = 8'h20;
    ff_ram[1949] = 8'h24;
    ff_ram[1950] = 8'h18;
    ff_ram[1951] = 8'h00;
    ff_ram[1952] = 8'h48;
    ff_ram[1953] = 8'h5C;
    ff_ram[1954] = 8'h6A;
    ff_ram[1955] = 8'hE2;
    ff_ram[1956] = 8'h24;
    ff_ram[1957] = 8'h10;
    ff_ram[1958] = 8'h10;
    ff_ram[1959] = 8'h00;
    ff_ram[1960] = 8'h10;
    ff_ram[1961] = 8'h9C;
    ff_ram[1962] = 8'hB2;
    ff_ram[1963] = 8'hD2;
    ff_ram[1964] = 8'h92;
    ff_ram[1965] = 8'h1C;
    ff_ram[1966] = 8'h20;
    ff_ram[1967] = 8'h00;
    ff_ram[1968] = 8'h10;
    ff_ram[1969] = 8'h1C;
    ff_ram[1970] = 8'h10;
    ff_ram[1971] = 8'h10;
    ff_ram[1972] = 8'h78;
    ff_ram[1973] = 8'h94;
    ff_ram[1974] = 8'h70;
    ff_ram[1975] = 8'h00;
    ff_ram[1976] = 8'h60;
    ff_ram[1977] = 8'h10;
    ff_ram[1978] = 8'h80;
    ff_ram[1979] = 8'hB8;
    ff_ram[1980] = 8'hC4;
    ff_ram[1981] = 8'h84;
    ff_ram[1982] = 8'h38;
    ff_ram[1983] = 8'h00;
    ff_ram[1984] = 8'h08;
    ff_ram[1985] = 8'h84;
    ff_ram[1986] = 8'h84;
    ff_ram[1987] = 8'h84;
    ff_ram[1988] = 8'h44;
    ff_ram[1989] = 8'h08;
    ff_ram[1990] = 8'h30;
    ff_ram[1991] = 8'h00;
    ff_ram[1992] = 8'h78;
    ff_ram[1993] = 8'h10;
    ff_ram[1994] = 8'h38;
    ff_ram[1995] = 8'h44;
    ff_ram[1996] = 8'hB4;
    ff_ram[1997] = 8'h4C;
    ff_ram[1998] = 8'h38;
    ff_ram[1999] = 8'h00;
    ff_ram[2000] = 8'h20;
    ff_ram[2001] = 8'h2C;
    ff_ram[2002] = 8'hF4;
    ff_ram[2003] = 8'h24;
    ff_ram[2004] = 8'h64;
    ff_ram[2005] = 8'hA4;
    ff_ram[2006] = 8'h26;
    ff_ram[2007] = 8'h00;
    ff_ram[2008] = 8'h78;
    ff_ram[2009] = 8'h10;
    ff_ram[2010] = 8'h20;
    ff_ram[2011] = 8'h78;
    ff_ram[2012] = 8'h84;
    ff_ram[2013] = 8'h04;
    ff_ram[2014] = 8'h38;
    ff_ram[2015] = 8'h00;
    ff_ram[2016] = 8'h40;
    ff_ram[2017] = 8'h40;
    ff_ram[2018] = 8'hDC;
    ff_ram[2019] = 8'h62;
    ff_ram[2020] = 8'h42;
    ff_ram[2021] = 8'hC2;
    ff_ram[2022] = 8'h44;
    ff_ram[2023] = 8'h00;
    ff_ram[2024] = 8'h10;
    ff_ram[2025] = 8'h10;
    ff_ram[2026] = 8'h20;
    ff_ram[2027] = 8'h20;
    ff_ram[2028] = 8'h60;
    ff_ram[2029] = 8'h52;
    ff_ram[2030] = 8'h8C;
    ff_ram[2031] = 8'h00;
    ff_ram[2032] = 8'h00;
    ff_ram[2033] = 8'h00;
    ff_ram[2034] = 8'h00;
    ff_ram[2035] = 8'h00;
    ff_ram[2036] = 8'h00;
    ff_ram[2037] = 8'h00;
    ff_ram[2038] = 8'h00;
    ff_ram[2039] = 8'h00;
    ff_ram[2040] = 8'hFF;
    ff_ram[2041] = 8'hFF;
    ff_ram[2042] = 8'hFF;
    ff_ram[2043] = 8'hFF;
    ff_ram[2044] = 8'hFF;
    ff_ram[2045] = 8'hFF;
    ff_ram[2046] = 8'hFF;
    ff_ram[2047] = 8'hFF;
    ff_ram[2048] = 8'h00;
    ff_ram[2049] = 8'h00;
    ff_ram[2050] = 8'h00;
    ff_ram[2051] = 8'h00;
    ff_ram[2052] = 8'h00;
    ff_ram[2053] = 8'h00;
    ff_ram[2054] = 8'h00;
    ff_ram[2055] = 8'h00;
    ff_ram[2056] = 8'h00;
    ff_ram[2057] = 8'h00;
    ff_ram[2058] = 8'h00;
    ff_ram[2059] = 8'h00;
    ff_ram[2060] = 8'h00;
    ff_ram[2061] = 8'h00;
    ff_ram[2062] = 8'h00;
    ff_ram[2063] = 8'h00;
    ff_ram[2064] = 8'h00;
    ff_ram[2065] = 8'h00;
    ff_ram[2066] = 8'h00;
    ff_ram[2067] = 8'h00;
    ff_ram[2068] = 8'h00;
    ff_ram[2069] = 8'h00;
    ff_ram[2070] = 8'h00;
    ff_ram[2071] = 8'h00;
    ff_ram[2072] = 8'h00;
    ff_ram[2073] = 8'h00;
    ff_ram[2074] = 8'h00;
    ff_ram[2075] = 8'h00;
    ff_ram[2076] = 8'h00;
    ff_ram[2077] = 8'h00;
    ff_ram[2078] = 8'h00;
    ff_ram[2079] = 8'h00;
    ff_ram[2080] = 8'h00;
    ff_ram[2081] = 8'h00;
    ff_ram[2082] = 8'h00;
    ff_ram[2083] = 8'h00;
    ff_ram[2084] = 8'h00;
    ff_ram[2085] = 8'h00;
    ff_ram[2086] = 8'h00;
    ff_ram[2087] = 8'h00;
    ff_ram[2088] = 8'h00;
    ff_ram[2089] = 8'h00;
    ff_ram[2090] = 8'h00;
    ff_ram[2091] = 8'h00;
    ff_ram[2092] = 8'h00;
    ff_ram[2093] = 8'h00;
    ff_ram[2094] = 8'h00;
    ff_ram[2095] = 8'h00;
    ff_ram[2096] = 8'h00;
    ff_ram[2097] = 8'h00;
    ff_ram[2098] = 8'h00;
    ff_ram[2099] = 8'h00;
    ff_ram[2100] = 8'h00;
    ff_ram[2101] = 8'h00;
    ff_ram[2102] = 8'h00;
    ff_ram[2103] = 8'h00;
    ff_ram[2104] = 8'h00;
    ff_ram[2105] = 8'h00;
    ff_ram[2106] = 8'h00;
    ff_ram[2107] = 8'h00;
    ff_ram[2108] = 8'h00;
    ff_ram[2109] = 8'h00;
    ff_ram[2110] = 8'h00;
    ff_ram[2111] = 8'h00;
    ff_ram[2112] = 8'h00;
    ff_ram[2113] = 8'h00;
    ff_ram[2114] = 8'h00;
    ff_ram[2115] = 8'h00;
    ff_ram[2116] = 8'h00;
    ff_ram[2117] = 8'h00;
    ff_ram[2118] = 8'h00;
    ff_ram[2119] = 8'h00;
    ff_ram[2120] = 8'h00;
    ff_ram[2121] = 8'h00;
    ff_ram[2122] = 8'h00;
    ff_ram[2123] = 8'h00;
    ff_ram[2124] = 8'h00;
    ff_ram[2125] = 8'h00;
    ff_ram[2126] = 8'h00;
    ff_ram[2127] = 8'h00;
    ff_ram[2128] = 8'h00;
    ff_ram[2129] = 8'h00;
    ff_ram[2130] = 8'h00;
    ff_ram[2131] = 8'h00;
    ff_ram[2132] = 8'h00;
    ff_ram[2133] = 8'h00;
    ff_ram[2134] = 8'h00;
    ff_ram[2135] = 8'h00;
    ff_ram[2136] = 8'h00;
    ff_ram[2137] = 8'h00;
    ff_ram[2138] = 8'h00;
    ff_ram[2139] = 8'h00;
    ff_ram[2140] = 8'h00;
    ff_ram[2141] = 8'h00;
    ff_ram[2142] = 8'h00;
    ff_ram[2143] = 8'h00;
    ff_ram[2144] = 8'h00;
    ff_ram[2145] = 8'h00;
    ff_ram[2146] = 8'h00;
    ff_ram[2147] = 8'h00;
    ff_ram[2148] = 8'h00;
    ff_ram[2149] = 8'h00;
    ff_ram[2150] = 8'h00;
    ff_ram[2151] = 8'h00;
    ff_ram[2152] = 8'h00;
    ff_ram[2153] = 8'h00;
    ff_ram[2154] = 8'h00;
    ff_ram[2155] = 8'h00;
    ff_ram[2156] = 8'h00;
    ff_ram[2157] = 8'h00;
    ff_ram[2158] = 8'h00;
    ff_ram[2159] = 8'h00;
    ff_ram[2160] = 8'h00;
    ff_ram[2161] = 8'h00;
    ff_ram[2162] = 8'h00;
    ff_ram[2163] = 8'h00;
    ff_ram[2164] = 8'h00;
    ff_ram[2165] = 8'h00;
    ff_ram[2166] = 8'h00;
    ff_ram[2167] = 8'h00;
    ff_ram[2168] = 8'h00;
    ff_ram[2169] = 8'h00;
    ff_ram[2170] = 8'h00;
    ff_ram[2171] = 8'h00;
    ff_ram[2172] = 8'h00;
    ff_ram[2173] = 8'h00;
    ff_ram[2174] = 8'h00;
    ff_ram[2175] = 8'h00;
    ff_ram[2176] = 8'h00;
    ff_ram[2177] = 8'h00;
    ff_ram[2178] = 8'h00;
    ff_ram[2179] = 8'h00;
    ff_ram[2180] = 8'h00;
    ff_ram[2181] = 8'h00;
    ff_ram[2182] = 8'h00;
    ff_ram[2183] = 8'h00;
    ff_ram[2184] = 8'h00;
    ff_ram[2185] = 8'h00;
    ff_ram[2186] = 8'h00;
    ff_ram[2187] = 8'h00;
    ff_ram[2188] = 8'h00;
    ff_ram[2189] = 8'h00;
    ff_ram[2190] = 8'h00;
    ff_ram[2191] = 8'h00;
    ff_ram[2192] = 8'h00;
    ff_ram[2193] = 8'h00;
    ff_ram[2194] = 8'h00;
    ff_ram[2195] = 8'h00;
    ff_ram[2196] = 8'h00;
    ff_ram[2197] = 8'h00;
    ff_ram[2198] = 8'h00;
    ff_ram[2199] = 8'h00;
    ff_ram[2200] = 8'h00;
    ff_ram[2201] = 8'h00;
    ff_ram[2202] = 8'h00;
    ff_ram[2203] = 8'h00;
    ff_ram[2204] = 8'h00;
    ff_ram[2205] = 8'h00;
    ff_ram[2206] = 8'h00;
    ff_ram[2207] = 8'h00;
    ff_ram[2208] = 8'h00;
    ff_ram[2209] = 8'h00;
    ff_ram[2210] = 8'h00;
    ff_ram[2211] = 8'h00;
    ff_ram[2212] = 8'h00;
    ff_ram[2213] = 8'h00;
    ff_ram[2214] = 8'h00;
    ff_ram[2215] = 8'h00;
    ff_ram[2216] = 8'h00;
    ff_ram[2217] = 8'h00;
    ff_ram[2218] = 8'h00;
    ff_ram[2219] = 8'h00;
    ff_ram[2220] = 8'h00;
    ff_ram[2221] = 8'h00;
    ff_ram[2222] = 8'h00;
    ff_ram[2223] = 8'h00;
    ff_ram[2224] = 8'h00;
    ff_ram[2225] = 8'h00;
    ff_ram[2226] = 8'h00;
    ff_ram[2227] = 8'h00;
    ff_ram[2228] = 8'h00;
    ff_ram[2229] = 8'h00;
    ff_ram[2230] = 8'h00;
    ff_ram[2231] = 8'h00;
    ff_ram[2232] = 8'h00;
    ff_ram[2233] = 8'h00;
    ff_ram[2234] = 8'h00;
    ff_ram[2235] = 8'h00;
    ff_ram[2236] = 8'h00;
    ff_ram[2237] = 8'h00;
    ff_ram[2238] = 8'h00;
    ff_ram[2239] = 8'h00;
    ff_ram[2240] = 8'h00;
    ff_ram[2241] = 8'h00;
    ff_ram[2242] = 8'h00;
    ff_ram[2243] = 8'h00;
    ff_ram[2244] = 8'h00;
    ff_ram[2245] = 8'h00;
    ff_ram[2246] = 8'h00;
    ff_ram[2247] = 8'h00;
    ff_ram[2248] = 8'h00;
    ff_ram[2249] = 8'h00;
    ff_ram[2250] = 8'h00;
    ff_ram[2251] = 8'h00;
    ff_ram[2252] = 8'h00;
    ff_ram[2253] = 8'h00;
    ff_ram[2254] = 8'h00;
    ff_ram[2255] = 8'h00;
    ff_ram[2256] = 8'h00;
    ff_ram[2257] = 8'h00;
    ff_ram[2258] = 8'h00;
    ff_ram[2259] = 8'h00;
    ff_ram[2260] = 8'h00;
    ff_ram[2261] = 8'h00;
    ff_ram[2262] = 8'h00;
    ff_ram[2263] = 8'h00;
    ff_ram[2264] = 8'h00;
    ff_ram[2265] = 8'h00;
    ff_ram[2266] = 8'h00;
    ff_ram[2267] = 8'h00;
    ff_ram[2268] = 8'h00;
    ff_ram[2269] = 8'h00;
    ff_ram[2270] = 8'h00;
    ff_ram[2271] = 8'h00;
    ff_ram[2272] = 8'h00;
    ff_ram[2273] = 8'h00;
    ff_ram[2274] = 8'h00;
    ff_ram[2275] = 8'h00;
    ff_ram[2276] = 8'h00;
    ff_ram[2277] = 8'h00;
    ff_ram[2278] = 8'h00;
    ff_ram[2279] = 8'h00;
    ff_ram[2280] = 8'h00;
    ff_ram[2281] = 8'h00;
    ff_ram[2282] = 8'h00;
    ff_ram[2283] = 8'h00;
    ff_ram[2284] = 8'h00;
    ff_ram[2285] = 8'h00;
    ff_ram[2286] = 8'h00;
    ff_ram[2287] = 8'h00;
    ff_ram[2288] = 8'h00;
    ff_ram[2289] = 8'h00;
    ff_ram[2290] = 8'h00;
    ff_ram[2291] = 8'h00;
    ff_ram[2292] = 8'h00;
    ff_ram[2293] = 8'h00;
    ff_ram[2294] = 8'h00;
    ff_ram[2295] = 8'h00;
    ff_ram[2296] = 8'h00;
    ff_ram[2297] = 8'h00;
    ff_ram[2298] = 8'h00;
    ff_ram[2299] = 8'h00;
    ff_ram[2300] = 8'h00;
    ff_ram[2301] = 8'h00;
    ff_ram[2302] = 8'h00;
    ff_ram[2303] = 8'h00;
    ff_ram[2304] = 8'h00;
    ff_ram[2305] = 8'h00;
    ff_ram[2306] = 8'h00;
    ff_ram[2307] = 8'h00;
    ff_ram[2308] = 8'h00;
    ff_ram[2309] = 8'h00;
    ff_ram[2310] = 8'h00;
    ff_ram[2311] = 8'h00;
    ff_ram[2312] = 8'h00;
    ff_ram[2313] = 8'h00;
    ff_ram[2314] = 8'h00;
    ff_ram[2315] = 8'h00;
    ff_ram[2316] = 8'h00;
    ff_ram[2317] = 8'h00;
    ff_ram[2318] = 8'h00;
    ff_ram[2319] = 8'h00;
    ff_ram[2320] = 8'h00;
    ff_ram[2321] = 8'h00;
    ff_ram[2322] = 8'h00;
    ff_ram[2323] = 8'h00;
    ff_ram[2324] = 8'h00;
    ff_ram[2325] = 8'h00;
    ff_ram[2326] = 8'h00;
    ff_ram[2327] = 8'h00;
    ff_ram[2328] = 8'h00;
    ff_ram[2329] = 8'h00;
    ff_ram[2330] = 8'h00;
    ff_ram[2331] = 8'h00;
    ff_ram[2332] = 8'h00;
    ff_ram[2333] = 8'h00;
    ff_ram[2334] = 8'h00;
    ff_ram[2335] = 8'h00;
    ff_ram[2336] = 8'h00;
    ff_ram[2337] = 8'h00;
    ff_ram[2338] = 8'h00;
    ff_ram[2339] = 8'h00;
    ff_ram[2340] = 8'h00;
    ff_ram[2341] = 8'h00;
    ff_ram[2342] = 8'h00;
    ff_ram[2343] = 8'h00;
    ff_ram[2344] = 8'h00;
    ff_ram[2345] = 8'h00;
    ff_ram[2346] = 8'h00;
    ff_ram[2347] = 8'h00;
    ff_ram[2348] = 8'h00;
    ff_ram[2349] = 8'h00;
    ff_ram[2350] = 8'h00;
    ff_ram[2351] = 8'h00;
    ff_ram[2352] = 8'h00;
    ff_ram[2353] = 8'h00;
    ff_ram[2354] = 8'h00;
    ff_ram[2355] = 8'h00;
    ff_ram[2356] = 8'h00;
    ff_ram[2357] = 8'h00;
    ff_ram[2358] = 8'h00;
    ff_ram[2359] = 8'h00;
    ff_ram[2360] = 8'h00;
    ff_ram[2361] = 8'h00;
    ff_ram[2362] = 8'h00;
    ff_ram[2363] = 8'h00;
    ff_ram[2364] = 8'h00;
    ff_ram[2365] = 8'h00;
    ff_ram[2366] = 8'h00;
    ff_ram[2367] = 8'h00;
    ff_ram[2368] = 8'h00;
    ff_ram[2369] = 8'h00;
    ff_ram[2370] = 8'h00;
    ff_ram[2371] = 8'h00;
    ff_ram[2372] = 8'h00;
    ff_ram[2373] = 8'h00;
    ff_ram[2374] = 8'h00;
    ff_ram[2375] = 8'h00;
    ff_ram[2376] = 8'h00;
    ff_ram[2377] = 8'h00;
    ff_ram[2378] = 8'h00;
    ff_ram[2379] = 8'h00;
    ff_ram[2380] = 8'h00;
    ff_ram[2381] = 8'h00;
    ff_ram[2382] = 8'h00;
    ff_ram[2383] = 8'h00;
    ff_ram[2384] = 8'h00;
    ff_ram[2385] = 8'h00;
    ff_ram[2386] = 8'h00;
    ff_ram[2387] = 8'h00;
    ff_ram[2388] = 8'h00;
    ff_ram[2389] = 8'h00;
    ff_ram[2390] = 8'h00;
    ff_ram[2391] = 8'h00;
    ff_ram[2392] = 8'h00;
    ff_ram[2393] = 8'h00;
    ff_ram[2394] = 8'h00;
    ff_ram[2395] = 8'h00;
    ff_ram[2396] = 8'h00;
    ff_ram[2397] = 8'h00;
    ff_ram[2398] = 8'h00;
    ff_ram[2399] = 8'h00;
    ff_ram[2400] = 8'h00;
    ff_ram[2401] = 8'h00;
    ff_ram[2402] = 8'h00;
    ff_ram[2403] = 8'h00;
    ff_ram[2404] = 8'h00;
    ff_ram[2405] = 8'h00;
    ff_ram[2406] = 8'h00;
    ff_ram[2407] = 8'h00;
    ff_ram[2408] = 8'h00;
    ff_ram[2409] = 8'h00;
    ff_ram[2410] = 8'h00;
    ff_ram[2411] = 8'h00;
    ff_ram[2412] = 8'h00;
    ff_ram[2413] = 8'h00;
    ff_ram[2414] = 8'h00;
    ff_ram[2415] = 8'h00;
    ff_ram[2416] = 8'h00;
    ff_ram[2417] = 8'h00;
    ff_ram[2418] = 8'h00;
    ff_ram[2419] = 8'h00;
    ff_ram[2420] = 8'h00;
    ff_ram[2421] = 8'h00;
    ff_ram[2422] = 8'h00;
    ff_ram[2423] = 8'h00;
    ff_ram[2424] = 8'h00;
    ff_ram[2425] = 8'h00;
    ff_ram[2426] = 8'h00;
    ff_ram[2427] = 8'h00;
    ff_ram[2428] = 8'h00;
    ff_ram[2429] = 8'h00;
    ff_ram[2430] = 8'h00;
    ff_ram[2431] = 8'h00;
    ff_ram[2432] = 8'h00;
    ff_ram[2433] = 8'h00;
    ff_ram[2434] = 8'h00;
    ff_ram[2435] = 8'h00;
    ff_ram[2436] = 8'h00;
    ff_ram[2437] = 8'h00;
    ff_ram[2438] = 8'h00;
    ff_ram[2439] = 8'h00;
    ff_ram[2440] = 8'h00;
    ff_ram[2441] = 8'h00;
    ff_ram[2442] = 8'h00;
    ff_ram[2443] = 8'h00;
    ff_ram[2444] = 8'h00;
    ff_ram[2445] = 8'h00;
    ff_ram[2446] = 8'h00;
    ff_ram[2447] = 8'h00;
    ff_ram[2448] = 8'h00;
    ff_ram[2449] = 8'h00;
    ff_ram[2450] = 8'h00;
    ff_ram[2451] = 8'h00;
    ff_ram[2452] = 8'h00;
    ff_ram[2453] = 8'h00;
    ff_ram[2454] = 8'h00;
    ff_ram[2455] = 8'h00;
    ff_ram[2456] = 8'h00;
    ff_ram[2457] = 8'h00;
    ff_ram[2458] = 8'h00;
    ff_ram[2459] = 8'h00;
    ff_ram[2460] = 8'h00;
    ff_ram[2461] = 8'h00;
    ff_ram[2462] = 8'h00;
    ff_ram[2463] = 8'h00;
    ff_ram[2464] = 8'h00;
    ff_ram[2465] = 8'h00;
    ff_ram[2466] = 8'h00;
    ff_ram[2467] = 8'h00;
    ff_ram[2468] = 8'h00;
    ff_ram[2469] = 8'h00;
    ff_ram[2470] = 8'h00;
    ff_ram[2471] = 8'h00;
    ff_ram[2472] = 8'h00;
    ff_ram[2473] = 8'h00;
    ff_ram[2474] = 8'h00;
    ff_ram[2475] = 8'h00;
    ff_ram[2476] = 8'h00;
    ff_ram[2477] = 8'h00;
    ff_ram[2478] = 8'h00;
    ff_ram[2479] = 8'h00;
    ff_ram[2480] = 8'h00;
    ff_ram[2481] = 8'h00;
    ff_ram[2482] = 8'h00;
    ff_ram[2483] = 8'h00;
    ff_ram[2484] = 8'h00;
    ff_ram[2485] = 8'h00;
    ff_ram[2486] = 8'h00;
    ff_ram[2487] = 8'h00;
    ff_ram[2488] = 8'h00;
    ff_ram[2489] = 8'h00;
    ff_ram[2490] = 8'h00;
    ff_ram[2491] = 8'h00;
    ff_ram[2492] = 8'h00;
    ff_ram[2493] = 8'h00;
    ff_ram[2494] = 8'h00;
    ff_ram[2495] = 8'h00;
    ff_ram[2496] = 8'h00;
    ff_ram[2497] = 8'h00;
    ff_ram[2498] = 8'h00;
    ff_ram[2499] = 8'h00;
    ff_ram[2500] = 8'h00;
    ff_ram[2501] = 8'h00;
    ff_ram[2502] = 8'h00;
    ff_ram[2503] = 8'h00;
    ff_ram[2504] = 8'h00;
    ff_ram[2505] = 8'h00;
    ff_ram[2506] = 8'h00;
    ff_ram[2507] = 8'h00;
    ff_ram[2508] = 8'h00;
    ff_ram[2509] = 8'h00;
    ff_ram[2510] = 8'h00;
    ff_ram[2511] = 8'h00;
    ff_ram[2512] = 8'h00;
    ff_ram[2513] = 8'h00;
    ff_ram[2514] = 8'h00;
    ff_ram[2515] = 8'h00;
    ff_ram[2516] = 8'h00;
    ff_ram[2517] = 8'h00;
    ff_ram[2518] = 8'h00;
    ff_ram[2519] = 8'h00;
    ff_ram[2520] = 8'h00;
    ff_ram[2521] = 8'h00;
    ff_ram[2522] = 8'h00;
    ff_ram[2523] = 8'h00;
    ff_ram[2524] = 8'h00;
    ff_ram[2525] = 8'h00;
    ff_ram[2526] = 8'h00;
    ff_ram[2527] = 8'h00;
    ff_ram[2528] = 8'h00;
    ff_ram[2529] = 8'h00;
    ff_ram[2530] = 8'h00;
    ff_ram[2531] = 8'h00;
    ff_ram[2532] = 8'h00;
    ff_ram[2533] = 8'h00;
    ff_ram[2534] = 8'h00;
    ff_ram[2535] = 8'h00;
    ff_ram[2536] = 8'h00;
    ff_ram[2537] = 8'h00;
    ff_ram[2538] = 8'h00;
    ff_ram[2539] = 8'h00;
    ff_ram[2540] = 8'h00;
    ff_ram[2541] = 8'h00;
    ff_ram[2542] = 8'h00;
    ff_ram[2543] = 8'h00;
    ff_ram[2544] = 8'h00;
    ff_ram[2545] = 8'h00;
    ff_ram[2546] = 8'h00;
    ff_ram[2547] = 8'h00;
    ff_ram[2548] = 8'h00;
    ff_ram[2549] = 8'h00;
    ff_ram[2550] = 8'h00;
    ff_ram[2551] = 8'h00;
    ff_ram[2552] = 8'h00;
    ff_ram[2553] = 8'h00;
    ff_ram[2554] = 8'h00;
    ff_ram[2555] = 8'h00;
    ff_ram[2556] = 8'h00;
    ff_ram[2557] = 8'h00;
    ff_ram[2558] = 8'h00;
    ff_ram[2559] = 8'h00;
    ff_ram[2560] = 8'h00;
    ff_ram[2561] = 8'h00;
    ff_ram[2562] = 8'h00;
    ff_ram[2563] = 8'h00;
    ff_ram[2564] = 8'h00;
    ff_ram[2565] = 8'h00;
    ff_ram[2566] = 8'h00;
    ff_ram[2567] = 8'h00;
    ff_ram[2568] = 8'h00;
    ff_ram[2569] = 8'h00;
    ff_ram[2570] = 8'h00;
    ff_ram[2571] = 8'h00;
    ff_ram[2572] = 8'h00;
    ff_ram[2573] = 8'h00;
    ff_ram[2574] = 8'h00;
    ff_ram[2575] = 8'h00;
    ff_ram[2576] = 8'h00;
    ff_ram[2577] = 8'h00;
    ff_ram[2578] = 8'h00;
    ff_ram[2579] = 8'h00;
    ff_ram[2580] = 8'h00;
    ff_ram[2581] = 8'h00;
    ff_ram[2582] = 8'h00;
    ff_ram[2583] = 8'h00;
    ff_ram[2584] = 8'h00;
    ff_ram[2585] = 8'h00;
    ff_ram[2586] = 8'h00;
    ff_ram[2587] = 8'h00;
    ff_ram[2588] = 8'h00;
    ff_ram[2589] = 8'h00;
    ff_ram[2590] = 8'h00;
    ff_ram[2591] = 8'h00;
    ff_ram[2592] = 8'h00;
    ff_ram[2593] = 8'h00;
    ff_ram[2594] = 8'h00;
    ff_ram[2595] = 8'h00;
    ff_ram[2596] = 8'h00;
    ff_ram[2597] = 8'h00;
    ff_ram[2598] = 8'h00;
    ff_ram[2599] = 8'h00;
    ff_ram[2600] = 8'h00;
    ff_ram[2601] = 8'h00;
    ff_ram[2602] = 8'h00;
    ff_ram[2603] = 8'h00;
    ff_ram[2604] = 8'h00;
    ff_ram[2605] = 8'h00;
    ff_ram[2606] = 8'h00;
    ff_ram[2607] = 8'h00;
    ff_ram[2608] = 8'h00;
    ff_ram[2609] = 8'h00;
    ff_ram[2610] = 8'h00;
    ff_ram[2611] = 8'h00;
    ff_ram[2612] = 8'h00;
    ff_ram[2613] = 8'h00;
    ff_ram[2614] = 8'h00;
    ff_ram[2615] = 8'h00;
    ff_ram[2616] = 8'h00;
    ff_ram[2617] = 8'h00;
    ff_ram[2618] = 8'h00;
    ff_ram[2619] = 8'h00;
    ff_ram[2620] = 8'h00;
    ff_ram[2621] = 8'h00;
    ff_ram[2622] = 8'h00;
    ff_ram[2623] = 8'h00;
    ff_ram[2624] = 8'h00;
    ff_ram[2625] = 8'h00;
    ff_ram[2626] = 8'h00;
    ff_ram[2627] = 8'h00;
    ff_ram[2628] = 8'h00;
    ff_ram[2629] = 8'h00;
    ff_ram[2630] = 8'h00;
    ff_ram[2631] = 8'h00;
    ff_ram[2632] = 8'h00;
    ff_ram[2633] = 8'h00;
    ff_ram[2634] = 8'h00;
    ff_ram[2635] = 8'h00;
    ff_ram[2636] = 8'h00;
    ff_ram[2637] = 8'h00;
    ff_ram[2638] = 8'h00;
    ff_ram[2639] = 8'h00;
    ff_ram[2640] = 8'h00;
    ff_ram[2641] = 8'h00;
    ff_ram[2642] = 8'h00;
    ff_ram[2643] = 8'h00;
    ff_ram[2644] = 8'h00;
    ff_ram[2645] = 8'h00;
    ff_ram[2646] = 8'h00;
    ff_ram[2647] = 8'h00;
    ff_ram[2648] = 8'h00;
    ff_ram[2649] = 8'h00;
    ff_ram[2650] = 8'h00;
    ff_ram[2651] = 8'h00;
    ff_ram[2652] = 8'h00;
    ff_ram[2653] = 8'h00;
    ff_ram[2654] = 8'h00;
    ff_ram[2655] = 8'h00;
    ff_ram[2656] = 8'h00;
    ff_ram[2657] = 8'h00;
    ff_ram[2658] = 8'h00;
    ff_ram[2659] = 8'h00;
    ff_ram[2660] = 8'h00;
    ff_ram[2661] = 8'h00;
    ff_ram[2662] = 8'h00;
    ff_ram[2663] = 8'h00;
    ff_ram[2664] = 8'h00;
    ff_ram[2665] = 8'h00;
    ff_ram[2666] = 8'h00;
    ff_ram[2667] = 8'h00;
    ff_ram[2668] = 8'h00;
    ff_ram[2669] = 8'h00;
    ff_ram[2670] = 8'h00;
    ff_ram[2671] = 8'h00;
    ff_ram[2672] = 8'h00;
    ff_ram[2673] = 8'h00;
    ff_ram[2674] = 8'h00;
    ff_ram[2675] = 8'h00;
    ff_ram[2676] = 8'h00;
    ff_ram[2677] = 8'h00;
    ff_ram[2678] = 8'h00;
    ff_ram[2679] = 8'h00;
    ff_ram[2680] = 8'h00;
    ff_ram[2681] = 8'h00;
    ff_ram[2682] = 8'h00;
    ff_ram[2683] = 8'h00;
    ff_ram[2684] = 8'h00;
    ff_ram[2685] = 8'h00;
    ff_ram[2686] = 8'h00;
    ff_ram[2687] = 8'h00;
    ff_ram[2688] = 8'h00;
    ff_ram[2689] = 8'h00;
    ff_ram[2690] = 8'h00;
    ff_ram[2691] = 8'h00;
    ff_ram[2692] = 8'h00;
    ff_ram[2693] = 8'h00;
    ff_ram[2694] = 8'h00;
    ff_ram[2695] = 8'h00;
    ff_ram[2696] = 8'h00;
    ff_ram[2697] = 8'h00;
    ff_ram[2698] = 8'h00;
    ff_ram[2699] = 8'h00;
    ff_ram[2700] = 8'h00;
    ff_ram[2701] = 8'h00;
    ff_ram[2702] = 8'h00;
    ff_ram[2703] = 8'h00;
    ff_ram[2704] = 8'h00;
    ff_ram[2705] = 8'h00;
    ff_ram[2706] = 8'h00;
    ff_ram[2707] = 8'h00;
    ff_ram[2708] = 8'h00;
    ff_ram[2709] = 8'h00;
    ff_ram[2710] = 8'h00;
    ff_ram[2711] = 8'h00;
    ff_ram[2712] = 8'h00;
    ff_ram[2713] = 8'h00;
    ff_ram[2714] = 8'h00;
    ff_ram[2715] = 8'h00;
    ff_ram[2716] = 8'h00;
    ff_ram[2717] = 8'h00;
    ff_ram[2718] = 8'h00;
    ff_ram[2719] = 8'h00;
    ff_ram[2720] = 8'h00;
    ff_ram[2721] = 8'h00;
    ff_ram[2722] = 8'h00;
    ff_ram[2723] = 8'h00;
    ff_ram[2724] = 8'h00;
    ff_ram[2725] = 8'h00;
    ff_ram[2726] = 8'h00;
    ff_ram[2727] = 8'h00;
    ff_ram[2728] = 8'h00;
    ff_ram[2729] = 8'h00;
    ff_ram[2730] = 8'h00;
    ff_ram[2731] = 8'h00;
    ff_ram[2732] = 8'h00;
    ff_ram[2733] = 8'h00;
    ff_ram[2734] = 8'h00;
    ff_ram[2735] = 8'h00;
    ff_ram[2736] = 8'h00;
    ff_ram[2737] = 8'h00;
    ff_ram[2738] = 8'h00;
    ff_ram[2739] = 8'h00;
    ff_ram[2740] = 8'h00;
    ff_ram[2741] = 8'h00;
    ff_ram[2742] = 8'h00;
    ff_ram[2743] = 8'h00;
    ff_ram[2744] = 8'h00;
    ff_ram[2745] = 8'h00;
    ff_ram[2746] = 8'h00;
    ff_ram[2747] = 8'h00;
    ff_ram[2748] = 8'h00;
    ff_ram[2749] = 8'h00;
    ff_ram[2750] = 8'h00;
    ff_ram[2751] = 8'h00;
    ff_ram[2752] = 8'h00;
    ff_ram[2753] = 8'h00;
    ff_ram[2754] = 8'h00;
    ff_ram[2755] = 8'h00;
    ff_ram[2756] = 8'h00;
    ff_ram[2757] = 8'h00;
    ff_ram[2758] = 8'h00;
    ff_ram[2759] = 8'h00;
    ff_ram[2760] = 8'h00;
    ff_ram[2761] = 8'h00;
    ff_ram[2762] = 8'h00;
    ff_ram[2763] = 8'h00;
    ff_ram[2764] = 8'h00;
    ff_ram[2765] = 8'h00;
    ff_ram[2766] = 8'h00;
    ff_ram[2767] = 8'h00;
    ff_ram[2768] = 8'h00;
    ff_ram[2769] = 8'h00;
    ff_ram[2770] = 8'h00;
    ff_ram[2771] = 8'h00;
    ff_ram[2772] = 8'h00;
    ff_ram[2773] = 8'h00;
    ff_ram[2774] = 8'h00;
    ff_ram[2775] = 8'h00;
    ff_ram[2776] = 8'h00;
    ff_ram[2777] = 8'h00;
    ff_ram[2778] = 8'h00;
    ff_ram[2779] = 8'h00;
    ff_ram[2780] = 8'h00;
    ff_ram[2781] = 8'h00;
    ff_ram[2782] = 8'h00;
    ff_ram[2783] = 8'h00;
    ff_ram[2784] = 8'h00;
    ff_ram[2785] = 8'h00;
    ff_ram[2786] = 8'h00;
    ff_ram[2787] = 8'h00;
    ff_ram[2788] = 8'h00;
    ff_ram[2789] = 8'h00;
    ff_ram[2790] = 8'h00;
    ff_ram[2791] = 8'h00;
    ff_ram[2792] = 8'h00;
    ff_ram[2793] = 8'h00;
    ff_ram[2794] = 8'h00;
    ff_ram[2795] = 8'h00;
    ff_ram[2796] = 8'h00;
    ff_ram[2797] = 8'h00;
    ff_ram[2798] = 8'h00;
    ff_ram[2799] = 8'h00;
    ff_ram[2800] = 8'h00;
    ff_ram[2801] = 8'h00;
    ff_ram[2802] = 8'h00;
    ff_ram[2803] = 8'h00;
    ff_ram[2804] = 8'h00;
    ff_ram[2805] = 8'h00;
    ff_ram[2806] = 8'h00;
    ff_ram[2807] = 8'h00;
    ff_ram[2808] = 8'h00;
    ff_ram[2809] = 8'h00;
    ff_ram[2810] = 8'h00;
    ff_ram[2811] = 8'h00;
    ff_ram[2812] = 8'h00;
    ff_ram[2813] = 8'h00;
    ff_ram[2814] = 8'h00;
    ff_ram[2815] = 8'h00;
    ff_ram[2816] = 8'h00;
    ff_ram[2817] = 8'h00;
    ff_ram[2818] = 8'h00;
    ff_ram[2819] = 8'h00;
    ff_ram[2820] = 8'h00;
    ff_ram[2821] = 8'h00;
    ff_ram[2822] = 8'h00;
    ff_ram[2823] = 8'h00;
    ff_ram[2824] = 8'h00;
    ff_ram[2825] = 8'h00;
    ff_ram[2826] = 8'h00;
    ff_ram[2827] = 8'h00;
    ff_ram[2828] = 8'h00;
    ff_ram[2829] = 8'h00;
    ff_ram[2830] = 8'h00;
    ff_ram[2831] = 8'h00;
    ff_ram[2832] = 8'h00;
    ff_ram[2833] = 8'h00;
    ff_ram[2834] = 8'h00;
    ff_ram[2835] = 8'h00;
    ff_ram[2836] = 8'h00;
    ff_ram[2837] = 8'h00;
    ff_ram[2838] = 8'h00;
    ff_ram[2839] = 8'h00;
    ff_ram[2840] = 8'h00;
    ff_ram[2841] = 8'h00;
    ff_ram[2842] = 8'h00;
    ff_ram[2843] = 8'h00;
    ff_ram[2844] = 8'h00;
    ff_ram[2845] = 8'h00;
    ff_ram[2846] = 8'h00;
    ff_ram[2847] = 8'h00;
    ff_ram[2848] = 8'h00;
    ff_ram[2849] = 8'h00;
    ff_ram[2850] = 8'h00;
    ff_ram[2851] = 8'h00;
    ff_ram[2852] = 8'h00;
    ff_ram[2853] = 8'h00;
    ff_ram[2854] = 8'h00;
    ff_ram[2855] = 8'h00;
    ff_ram[2856] = 8'h00;
    ff_ram[2857] = 8'h00;
    ff_ram[2858] = 8'h00;
    ff_ram[2859] = 8'h00;
    ff_ram[2860] = 8'h00;
    ff_ram[2861] = 8'h00;
    ff_ram[2862] = 8'h00;
    ff_ram[2863] = 8'h00;
    ff_ram[2864] = 8'h00;
    ff_ram[2865] = 8'h00;
    ff_ram[2866] = 8'h00;
    ff_ram[2867] = 8'h00;
    ff_ram[2868] = 8'h00;
    ff_ram[2869] = 8'h00;
    ff_ram[2870] = 8'h00;
    ff_ram[2871] = 8'h00;
    ff_ram[2872] = 8'h00;
    ff_ram[2873] = 8'h00;
    ff_ram[2874] = 8'h00;
    ff_ram[2875] = 8'h00;
    ff_ram[2876] = 8'h00;
    ff_ram[2877] = 8'h00;
    ff_ram[2878] = 8'h00;
    ff_ram[2879] = 8'h00;
    ff_ram[2880] = 8'h00;
    ff_ram[2881] = 8'h00;
    ff_ram[2882] = 8'h00;
    ff_ram[2883] = 8'h00;
    ff_ram[2884] = 8'h00;
    ff_ram[2885] = 8'h00;
    ff_ram[2886] = 8'h00;
    ff_ram[2887] = 8'h00;
    ff_ram[2888] = 8'h00;
    ff_ram[2889] = 8'h00;
    ff_ram[2890] = 8'h00;
    ff_ram[2891] = 8'h00;
    ff_ram[2892] = 8'h00;
    ff_ram[2893] = 8'h00;
    ff_ram[2894] = 8'h00;
    ff_ram[2895] = 8'h00;
    ff_ram[2896] = 8'h00;
    ff_ram[2897] = 8'h00;
    ff_ram[2898] = 8'h00;
    ff_ram[2899] = 8'h00;
    ff_ram[2900] = 8'h00;
    ff_ram[2901] = 8'h00;
    ff_ram[2902] = 8'h00;
    ff_ram[2903] = 8'h00;
    ff_ram[2904] = 8'h00;
    ff_ram[2905] = 8'h00;
    ff_ram[2906] = 8'h00;
    ff_ram[2907] = 8'h00;
    ff_ram[2908] = 8'h00;
    ff_ram[2909] = 8'h00;
    ff_ram[2910] = 8'h00;
    ff_ram[2911] = 8'h00;
    ff_ram[2912] = 8'h00;
    ff_ram[2913] = 8'h00;
    ff_ram[2914] = 8'h00;
    ff_ram[2915] = 8'h00;
    ff_ram[2916] = 8'h00;
    ff_ram[2917] = 8'h00;
    ff_ram[2918] = 8'h00;
    ff_ram[2919] = 8'h00;
    ff_ram[2920] = 8'h00;
    ff_ram[2921] = 8'h00;
    ff_ram[2922] = 8'h00;
    ff_ram[2923] = 8'h00;
    ff_ram[2924] = 8'h00;
    ff_ram[2925] = 8'h00;
    ff_ram[2926] = 8'h00;
    ff_ram[2927] = 8'h00;
    ff_ram[2928] = 8'h00;
    ff_ram[2929] = 8'h00;
    ff_ram[2930] = 8'h00;
    ff_ram[2931] = 8'h00;
    ff_ram[2932] = 8'h00;
    ff_ram[2933] = 8'h00;
    ff_ram[2934] = 8'h00;
    ff_ram[2935] = 8'h00;
    ff_ram[2936] = 8'h00;
    ff_ram[2937] = 8'h00;
    ff_ram[2938] = 8'h00;
    ff_ram[2939] = 8'h00;
    ff_ram[2940] = 8'h00;
    ff_ram[2941] = 8'h00;
    ff_ram[2942] = 8'h00;
    ff_ram[2943] = 8'h00;
    ff_ram[2944] = 8'h00;
    ff_ram[2945] = 8'h00;
    ff_ram[2946] = 8'h00;
    ff_ram[2947] = 8'h00;
    ff_ram[2948] = 8'h00;
    ff_ram[2949] = 8'h00;
    ff_ram[2950] = 8'h00;
    ff_ram[2951] = 8'h00;
    ff_ram[2952] = 8'h00;
    ff_ram[2953] = 8'h00;
    ff_ram[2954] = 8'h00;
    ff_ram[2955] = 8'h00;
    ff_ram[2956] = 8'h00;
    ff_ram[2957] = 8'h00;
    ff_ram[2958] = 8'h00;
    ff_ram[2959] = 8'h00;
    ff_ram[2960] = 8'h00;
    ff_ram[2961] = 8'h00;
    ff_ram[2962] = 8'h00;
    ff_ram[2963] = 8'h00;
    ff_ram[2964] = 8'h00;
    ff_ram[2965] = 8'h00;
    ff_ram[2966] = 8'h00;
    ff_ram[2967] = 8'h00;
    ff_ram[2968] = 8'h00;
    ff_ram[2969] = 8'h00;
    ff_ram[2970] = 8'h00;
    ff_ram[2971] = 8'h00;
    ff_ram[2972] = 8'h00;
    ff_ram[2973] = 8'h00;
    ff_ram[2974] = 8'h00;
    ff_ram[2975] = 8'h00;
    ff_ram[2976] = 8'h00;
    ff_ram[2977] = 8'h00;
    ff_ram[2978] = 8'h00;
    ff_ram[2979] = 8'h00;
    ff_ram[2980] = 8'h00;
    ff_ram[2981] = 8'h00;
    ff_ram[2982] = 8'h00;
    ff_ram[2983] = 8'h00;
    ff_ram[2984] = 8'h00;
    ff_ram[2985] = 8'h00;
    ff_ram[2986] = 8'h00;
    ff_ram[2987] = 8'h00;
    ff_ram[2988] = 8'h00;
    ff_ram[2989] = 8'h00;
    ff_ram[2990] = 8'h00;
    ff_ram[2991] = 8'h00;
    ff_ram[2992] = 8'h00;
    ff_ram[2993] = 8'h00;
    ff_ram[2994] = 8'h00;
    ff_ram[2995] = 8'h00;
    ff_ram[2996] = 8'h00;
    ff_ram[2997] = 8'h00;
    ff_ram[2998] = 8'h00;
    ff_ram[2999] = 8'h00;
    ff_ram[3000] = 8'h00;
    ff_ram[3001] = 8'h00;
    ff_ram[3002] = 8'h00;
    ff_ram[3003] = 8'h00;
    ff_ram[3004] = 8'h00;
    ff_ram[3005] = 8'h00;
    ff_ram[3006] = 8'h00;
    ff_ram[3007] = 8'h00;
    ff_ram[3008] = 8'h00;
    ff_ram[3009] = 8'h00;
    ff_ram[3010] = 8'h00;
    ff_ram[3011] = 8'h00;
    ff_ram[3012] = 8'h00;
    ff_ram[3013] = 8'h00;
    ff_ram[3014] = 8'h00;
    ff_ram[3015] = 8'h00;
    ff_ram[3016] = 8'h00;
    ff_ram[3017] = 8'h00;
    ff_ram[3018] = 8'h00;
    ff_ram[3019] = 8'h00;
    ff_ram[3020] = 8'h00;
    ff_ram[3021] = 8'h00;
    ff_ram[3022] = 8'h00;
    ff_ram[3023] = 8'h00;
    ff_ram[3024] = 8'h00;
    ff_ram[3025] = 8'h00;
    ff_ram[3026] = 8'h00;
    ff_ram[3027] = 8'h00;
    ff_ram[3028] = 8'h00;
    ff_ram[3029] = 8'h00;
    ff_ram[3030] = 8'h00;
    ff_ram[3031] = 8'h00;
    ff_ram[3032] = 8'h00;
    ff_ram[3033] = 8'h00;
    ff_ram[3034] = 8'h00;
    ff_ram[3035] = 8'h00;
    ff_ram[3036] = 8'h00;
    ff_ram[3037] = 8'h00;
    ff_ram[3038] = 8'h00;
    ff_ram[3039] = 8'h00;
    ff_ram[3040] = 8'h00;
    ff_ram[3041] = 8'h00;
    ff_ram[3042] = 8'h00;
    ff_ram[3043] = 8'h00;
    ff_ram[3044] = 8'h00;
    ff_ram[3045] = 8'h00;
    ff_ram[3046] = 8'h00;
    ff_ram[3047] = 8'h00;
    ff_ram[3048] = 8'h00;
    ff_ram[3049] = 8'h00;
    ff_ram[3050] = 8'h00;
    ff_ram[3051] = 8'h00;
    ff_ram[3052] = 8'h00;
    ff_ram[3053] = 8'h00;
    ff_ram[3054] = 8'h00;
    ff_ram[3055] = 8'h00;
    ff_ram[3056] = 8'h00;
    ff_ram[3057] = 8'h00;
    ff_ram[3058] = 8'h00;
    ff_ram[3059] = 8'h00;
    ff_ram[3060] = 8'h00;
    ff_ram[3061] = 8'h00;
    ff_ram[3062] = 8'h00;
    ff_ram[3063] = 8'h00;
    ff_ram[3064] = 8'h00;
    ff_ram[3065] = 8'h00;
    ff_ram[3066] = 8'h00;
    ff_ram[3067] = 8'h00;
    ff_ram[3068] = 8'h00;
    ff_ram[3069] = 8'h00;
    ff_ram[3070] = 8'h00;
    ff_ram[3071] = 8'h00;
    ff_ram[3072] = 8'h00;
    ff_ram[3073] = 8'h00;
    ff_ram[3074] = 8'h00;
    ff_ram[3075] = 8'h00;
    ff_ram[3076] = 8'h00;
    ff_ram[3077] = 8'h00;
    ff_ram[3078] = 8'h00;
    ff_ram[3079] = 8'h00;
    ff_ram[3080] = 8'h00;
    ff_ram[3081] = 8'h00;
    ff_ram[3082] = 8'h00;
    ff_ram[3083] = 8'h00;
    ff_ram[3084] = 8'h00;
    ff_ram[3085] = 8'h00;
    ff_ram[3086] = 8'h00;
    ff_ram[3087] = 8'h00;
    ff_ram[3088] = 8'h00;
    ff_ram[3089] = 8'h00;
    ff_ram[3090] = 8'h00;
    ff_ram[3091] = 8'h00;
    ff_ram[3092] = 8'h00;
    ff_ram[3093] = 8'h00;
    ff_ram[3094] = 8'h00;
    ff_ram[3095] = 8'h00;
    ff_ram[3096] = 8'h00;
    ff_ram[3097] = 8'h00;
    ff_ram[3098] = 8'h00;
    ff_ram[3099] = 8'h00;
    ff_ram[3100] = 8'h00;
    ff_ram[3101] = 8'h00;
    ff_ram[3102] = 8'h00;
    ff_ram[3103] = 8'h00;
    ff_ram[3104] = 8'h00;
    ff_ram[3105] = 8'h00;
    ff_ram[3106] = 8'h00;
    ff_ram[3107] = 8'h00;
    ff_ram[3108] = 8'h00;
    ff_ram[3109] = 8'h00;
    ff_ram[3110] = 8'h00;
    ff_ram[3111] = 8'h00;
    ff_ram[3112] = 8'h00;
    ff_ram[3113] = 8'h00;
    ff_ram[3114] = 8'h00;
    ff_ram[3115] = 8'h00;
    ff_ram[3116] = 8'h00;
    ff_ram[3117] = 8'h00;
    ff_ram[3118] = 8'h00;
    ff_ram[3119] = 8'h00;
    ff_ram[3120] = 8'h00;
    ff_ram[3121] = 8'h00;
    ff_ram[3122] = 8'h00;
    ff_ram[3123] = 8'h00;
    ff_ram[3124] = 8'h00;
    ff_ram[3125] = 8'h00;
    ff_ram[3126] = 8'h00;
    ff_ram[3127] = 8'h00;
    ff_ram[3128] = 8'h00;
    ff_ram[3129] = 8'h00;
    ff_ram[3130] = 8'h00;
    ff_ram[3131] = 8'h00;
    ff_ram[3132] = 8'h00;
    ff_ram[3133] = 8'h00;
    ff_ram[3134] = 8'h00;
    ff_ram[3135] = 8'h00;
    ff_ram[3136] = 8'h00;
    ff_ram[3137] = 8'h00;
    ff_ram[3138] = 8'h00;
    ff_ram[3139] = 8'h00;
    ff_ram[3140] = 8'h00;
    ff_ram[3141] = 8'h00;
    ff_ram[3142] = 8'h00;
    ff_ram[3143] = 8'h00;
    ff_ram[3144] = 8'h00;
    ff_ram[3145] = 8'h00;
    ff_ram[3146] = 8'h00;
    ff_ram[3147] = 8'h00;
    ff_ram[3148] = 8'h00;
    ff_ram[3149] = 8'h00;
    ff_ram[3150] = 8'h00;
    ff_ram[3151] = 8'h00;
    ff_ram[3152] = 8'h00;
    ff_ram[3153] = 8'h00;
    ff_ram[3154] = 8'h00;
    ff_ram[3155] = 8'h00;
    ff_ram[3156] = 8'h00;
    ff_ram[3157] = 8'h00;
    ff_ram[3158] = 8'h00;
    ff_ram[3159] = 8'h00;
    ff_ram[3160] = 8'h00;
    ff_ram[3161] = 8'h00;
    ff_ram[3162] = 8'h00;
    ff_ram[3163] = 8'h00;
    ff_ram[3164] = 8'h00;
    ff_ram[3165] = 8'h00;
    ff_ram[3166] = 8'h00;
    ff_ram[3167] = 8'h00;
    ff_ram[3168] = 8'h00;
    ff_ram[3169] = 8'h00;
    ff_ram[3170] = 8'h00;
    ff_ram[3171] = 8'h00;
    ff_ram[3172] = 8'h00;
    ff_ram[3173] = 8'h00;
    ff_ram[3174] = 8'h00;
    ff_ram[3175] = 8'h00;
    ff_ram[3176] = 8'h00;
    ff_ram[3177] = 8'h00;
    ff_ram[3178] = 8'h00;
    ff_ram[3179] = 8'h00;
    ff_ram[3180] = 8'h00;
    ff_ram[3181] = 8'h00;
    ff_ram[3182] = 8'h00;
    ff_ram[3183] = 8'h00;
    ff_ram[3184] = 8'h00;
    ff_ram[3185] = 8'h00;
    ff_ram[3186] = 8'h00;
    ff_ram[3187] = 8'h00;
    ff_ram[3188] = 8'h00;
    ff_ram[3189] = 8'h00;
    ff_ram[3190] = 8'h00;
    ff_ram[3191] = 8'h00;
    ff_ram[3192] = 8'h00;
    ff_ram[3193] = 8'h00;
    ff_ram[3194] = 8'h00;
    ff_ram[3195] = 8'h00;
    ff_ram[3196] = 8'h00;
    ff_ram[3197] = 8'h00;
    ff_ram[3198] = 8'h00;
    ff_ram[3199] = 8'h00;
    ff_ram[3200] = 8'h00;
    ff_ram[3201] = 8'h00;
    ff_ram[3202] = 8'h00;
    ff_ram[3203] = 8'h00;
    ff_ram[3204] = 8'h00;
    ff_ram[3205] = 8'h00;
    ff_ram[3206] = 8'h00;
    ff_ram[3207] = 8'h00;
    ff_ram[3208] = 8'h00;
    ff_ram[3209] = 8'h00;
    ff_ram[3210] = 8'h00;
    ff_ram[3211] = 8'h00;
    ff_ram[3212] = 8'h00;
    ff_ram[3213] = 8'h00;
    ff_ram[3214] = 8'h00;
    ff_ram[3215] = 8'h00;
    ff_ram[3216] = 8'h00;
    ff_ram[3217] = 8'h00;
    ff_ram[3218] = 8'h00;
    ff_ram[3219] = 8'h00;
    ff_ram[3220] = 8'h00;
    ff_ram[3221] = 8'h00;
    ff_ram[3222] = 8'h00;
    ff_ram[3223] = 8'h00;
    ff_ram[3224] = 8'h00;
    ff_ram[3225] = 8'h00;
    ff_ram[3226] = 8'h00;
    ff_ram[3227] = 8'h00;
    ff_ram[3228] = 8'h00;
    ff_ram[3229] = 8'h00;
    ff_ram[3230] = 8'h00;
    ff_ram[3231] = 8'h00;
    ff_ram[3232] = 8'h00;
    ff_ram[3233] = 8'h00;
    ff_ram[3234] = 8'h00;
    ff_ram[3235] = 8'h00;
    ff_ram[3236] = 8'h00;
    ff_ram[3237] = 8'h00;
    ff_ram[3238] = 8'h00;
    ff_ram[3239] = 8'h00;
    ff_ram[3240] = 8'h00;
    ff_ram[3241] = 8'h00;
    ff_ram[3242] = 8'h00;
    ff_ram[3243] = 8'h00;
    ff_ram[3244] = 8'h00;
    ff_ram[3245] = 8'h00;
    ff_ram[3246] = 8'h00;
    ff_ram[3247] = 8'h00;
    ff_ram[3248] = 8'h00;
    ff_ram[3249] = 8'h00;
    ff_ram[3250] = 8'h00;
    ff_ram[3251] = 8'h00;
    ff_ram[3252] = 8'h00;
    ff_ram[3253] = 8'h00;
    ff_ram[3254] = 8'h00;
    ff_ram[3255] = 8'h00;
    ff_ram[3256] = 8'h00;
    ff_ram[3257] = 8'h00;
    ff_ram[3258] = 8'h00;
    ff_ram[3259] = 8'h00;
    ff_ram[3260] = 8'h00;
    ff_ram[3261] = 8'h00;
    ff_ram[3262] = 8'h00;
    ff_ram[3263] = 8'h00;
    ff_ram[3264] = 8'h00;
    ff_ram[3265] = 8'h00;
    ff_ram[3266] = 8'h00;
    ff_ram[3267] = 8'h00;
    ff_ram[3268] = 8'h00;
    ff_ram[3269] = 8'h00;
    ff_ram[3270] = 8'h00;
    ff_ram[3271] = 8'h00;
    ff_ram[3272] = 8'h00;
    ff_ram[3273] = 8'h00;
    ff_ram[3274] = 8'h00;
    ff_ram[3275] = 8'h00;
    ff_ram[3276] = 8'h00;
    ff_ram[3277] = 8'h00;
    ff_ram[3278] = 8'h00;
    ff_ram[3279] = 8'h00;
    ff_ram[3280] = 8'h00;
    ff_ram[3281] = 8'h00;
    ff_ram[3282] = 8'h00;
    ff_ram[3283] = 8'h00;
    ff_ram[3284] = 8'h00;
    ff_ram[3285] = 8'h00;
    ff_ram[3286] = 8'h00;
    ff_ram[3287] = 8'h00;
    ff_ram[3288] = 8'h00;
    ff_ram[3289] = 8'h00;
    ff_ram[3290] = 8'h00;
    ff_ram[3291] = 8'h00;
    ff_ram[3292] = 8'h00;
    ff_ram[3293] = 8'h00;
    ff_ram[3294] = 8'h00;
    ff_ram[3295] = 8'h00;
    ff_ram[3296] = 8'h00;
    ff_ram[3297] = 8'h00;
    ff_ram[3298] = 8'h00;
    ff_ram[3299] = 8'h00;
    ff_ram[3300] = 8'h00;
    ff_ram[3301] = 8'h00;
    ff_ram[3302] = 8'h00;
    ff_ram[3303] = 8'h00;
    ff_ram[3304] = 8'h00;
    ff_ram[3305] = 8'h00;
    ff_ram[3306] = 8'h00;
    ff_ram[3307] = 8'h00;
    ff_ram[3308] = 8'h00;
    ff_ram[3309] = 8'h00;
    ff_ram[3310] = 8'h00;
    ff_ram[3311] = 8'h00;
    ff_ram[3312] = 8'h00;
    ff_ram[3313] = 8'h00;
    ff_ram[3314] = 8'h00;
    ff_ram[3315] = 8'h00;
    ff_ram[3316] = 8'h00;
    ff_ram[3317] = 8'h00;
    ff_ram[3318] = 8'h00;
    ff_ram[3319] = 8'h00;
    ff_ram[3320] = 8'h00;
    ff_ram[3321] = 8'h00;
    ff_ram[3322] = 8'h00;
    ff_ram[3323] = 8'h00;
    ff_ram[3324] = 8'h00;
    ff_ram[3325] = 8'h00;
    ff_ram[3326] = 8'h00;
    ff_ram[3327] = 8'h00;
    ff_ram[3328] = 8'h00;
    ff_ram[3329] = 8'h00;
    ff_ram[3330] = 8'h00;
    ff_ram[3331] = 8'h00;
    ff_ram[3332] = 8'h00;
    ff_ram[3333] = 8'h00;
    ff_ram[3334] = 8'h00;
    ff_ram[3335] = 8'h00;
    ff_ram[3336] = 8'h00;
    ff_ram[3337] = 8'h00;
    ff_ram[3338] = 8'h00;
    ff_ram[3339] = 8'h00;
    ff_ram[3340] = 8'h00;
    ff_ram[3341] = 8'h00;
    ff_ram[3342] = 8'h00;
    ff_ram[3343] = 8'h00;
    ff_ram[3344] = 8'h00;
    ff_ram[3345] = 8'h00;
    ff_ram[3346] = 8'h00;
    ff_ram[3347] = 8'h00;
    ff_ram[3348] = 8'h00;
    ff_ram[3349] = 8'h00;
    ff_ram[3350] = 8'h00;
    ff_ram[3351] = 8'h00;
    ff_ram[3352] = 8'h00;
    ff_ram[3353] = 8'h00;
    ff_ram[3354] = 8'h00;
    ff_ram[3355] = 8'h00;
    ff_ram[3356] = 8'h00;
    ff_ram[3357] = 8'h00;
    ff_ram[3358] = 8'h00;
    ff_ram[3359] = 8'h00;
    ff_ram[3360] = 8'h00;
    ff_ram[3361] = 8'h00;
    ff_ram[3362] = 8'h00;
    ff_ram[3363] = 8'h00;
    ff_ram[3364] = 8'h00;
    ff_ram[3365] = 8'h00;
    ff_ram[3366] = 8'h00;
    ff_ram[3367] = 8'h00;
    ff_ram[3368] = 8'h00;
    ff_ram[3369] = 8'h00;
    ff_ram[3370] = 8'h00;
    ff_ram[3371] = 8'h00;
    ff_ram[3372] = 8'h00;
    ff_ram[3373] = 8'h00;
    ff_ram[3374] = 8'h00;
    ff_ram[3375] = 8'h00;
    ff_ram[3376] = 8'h00;
    ff_ram[3377] = 8'h00;
    ff_ram[3378] = 8'h00;
    ff_ram[3379] = 8'h00;
    ff_ram[3380] = 8'h00;
    ff_ram[3381] = 8'h00;
    ff_ram[3382] = 8'h00;
    ff_ram[3383] = 8'h00;
    ff_ram[3384] = 8'h00;
    ff_ram[3385] = 8'h00;
    ff_ram[3386] = 8'h00;
    ff_ram[3387] = 8'h00;
    ff_ram[3388] = 8'h00;
    ff_ram[3389] = 8'h00;
    ff_ram[3390] = 8'h00;
    ff_ram[3391] = 8'h00;
    ff_ram[3392] = 8'h00;
    ff_ram[3393] = 8'h00;
    ff_ram[3394] = 8'h00;
    ff_ram[3395] = 8'h00;
    ff_ram[3396] = 8'h00;
    ff_ram[3397] = 8'h00;
    ff_ram[3398] = 8'h00;
    ff_ram[3399] = 8'h00;
    ff_ram[3400] = 8'h00;
    ff_ram[3401] = 8'h00;
    ff_ram[3402] = 8'h00;
    ff_ram[3403] = 8'h00;
    ff_ram[3404] = 8'h00;
    ff_ram[3405] = 8'h00;
    ff_ram[3406] = 8'h00;
    ff_ram[3407] = 8'h00;
    ff_ram[3408] = 8'h00;
    ff_ram[3409] = 8'h00;
    ff_ram[3410] = 8'h00;
    ff_ram[3411] = 8'h00;
    ff_ram[3412] = 8'h00;
    ff_ram[3413] = 8'h00;
    ff_ram[3414] = 8'h00;
    ff_ram[3415] = 8'h00;
    ff_ram[3416] = 8'h00;
    ff_ram[3417] = 8'h00;
    ff_ram[3418] = 8'h00;
    ff_ram[3419] = 8'h00;
    ff_ram[3420] = 8'h00;
    ff_ram[3421] = 8'h00;
    ff_ram[3422] = 8'h00;
    ff_ram[3423] = 8'h00;
    ff_ram[3424] = 8'h00;
    ff_ram[3425] = 8'h00;
    ff_ram[3426] = 8'h00;
    ff_ram[3427] = 8'h00;
    ff_ram[3428] = 8'h00;
    ff_ram[3429] = 8'h00;
    ff_ram[3430] = 8'h00;
    ff_ram[3431] = 8'h00;
    ff_ram[3432] = 8'h00;
    ff_ram[3433] = 8'h00;
    ff_ram[3434] = 8'h00;
    ff_ram[3435] = 8'h00;
    ff_ram[3436] = 8'h00;
    ff_ram[3437] = 8'h00;
    ff_ram[3438] = 8'h00;
    ff_ram[3439] = 8'h00;
    ff_ram[3440] = 8'h00;
    ff_ram[3441] = 8'h00;
    ff_ram[3442] = 8'h00;
    ff_ram[3443] = 8'h00;
    ff_ram[3444] = 8'h00;
    ff_ram[3445] = 8'h00;
    ff_ram[3446] = 8'h00;
    ff_ram[3447] = 8'h00;
    ff_ram[3448] = 8'h00;
    ff_ram[3449] = 8'h00;
    ff_ram[3450] = 8'h00;
    ff_ram[3451] = 8'h00;
    ff_ram[3452] = 8'h00;
    ff_ram[3453] = 8'h00;
    ff_ram[3454] = 8'h00;
    ff_ram[3455] = 8'h00;
    ff_ram[3456] = 8'h00;
    ff_ram[3457] = 8'h00;
    ff_ram[3458] = 8'h00;
    ff_ram[3459] = 8'h00;
    ff_ram[3460] = 8'h00;
    ff_ram[3461] = 8'h00;
    ff_ram[3462] = 8'h00;
    ff_ram[3463] = 8'h00;
    ff_ram[3464] = 8'h00;
    ff_ram[3465] = 8'h00;
    ff_ram[3466] = 8'h00;
    ff_ram[3467] = 8'h00;
    ff_ram[3468] = 8'h00;
    ff_ram[3469] = 8'h00;
    ff_ram[3470] = 8'h00;
    ff_ram[3471] = 8'h00;
    ff_ram[3472] = 8'h00;
    ff_ram[3473] = 8'h00;
    ff_ram[3474] = 8'h00;
    ff_ram[3475] = 8'h00;
    ff_ram[3476] = 8'h00;
    ff_ram[3477] = 8'h00;
    ff_ram[3478] = 8'h00;
    ff_ram[3479] = 8'h00;
    ff_ram[3480] = 8'h00;
    ff_ram[3481] = 8'h00;
    ff_ram[3482] = 8'h00;
    ff_ram[3483] = 8'h00;
    ff_ram[3484] = 8'h00;
    ff_ram[3485] = 8'h00;
    ff_ram[3486] = 8'h00;
    ff_ram[3487] = 8'h00;
    ff_ram[3488] = 8'h00;
    ff_ram[3489] = 8'h00;
    ff_ram[3490] = 8'h00;
    ff_ram[3491] = 8'h00;
    ff_ram[3492] = 8'h00;
    ff_ram[3493] = 8'h00;
    ff_ram[3494] = 8'h00;
    ff_ram[3495] = 8'h00;
    ff_ram[3496] = 8'h00;
    ff_ram[3497] = 8'h00;
    ff_ram[3498] = 8'h00;
    ff_ram[3499] = 8'h00;
    ff_ram[3500] = 8'h00;
    ff_ram[3501] = 8'h00;
    ff_ram[3502] = 8'h00;
    ff_ram[3503] = 8'h00;
    ff_ram[3504] = 8'h00;
    ff_ram[3505] = 8'h00;
    ff_ram[3506] = 8'h00;
    ff_ram[3507] = 8'h00;
    ff_ram[3508] = 8'h00;
    ff_ram[3509] = 8'h00;
    ff_ram[3510] = 8'h00;
    ff_ram[3511] = 8'h00;
    ff_ram[3512] = 8'h00;
    ff_ram[3513] = 8'h00;
    ff_ram[3514] = 8'h00;
    ff_ram[3515] = 8'h00;
    ff_ram[3516] = 8'h00;
    ff_ram[3517] = 8'h00;
    ff_ram[3518] = 8'h00;
    ff_ram[3519] = 8'h00;
    ff_ram[3520] = 8'h00;
    ff_ram[3521] = 8'h00;
    ff_ram[3522] = 8'h00;
    ff_ram[3523] = 8'h00;
    ff_ram[3524] = 8'h00;
    ff_ram[3525] = 8'h00;
    ff_ram[3526] = 8'h00;
    ff_ram[3527] = 8'h00;
    ff_ram[3528] = 8'h00;
    ff_ram[3529] = 8'h00;
    ff_ram[3530] = 8'h00;
    ff_ram[3531] = 8'h00;
    ff_ram[3532] = 8'h00;
    ff_ram[3533] = 8'h00;
    ff_ram[3534] = 8'h00;
    ff_ram[3535] = 8'h00;
    ff_ram[3536] = 8'h00;
    ff_ram[3537] = 8'h00;
    ff_ram[3538] = 8'h00;
    ff_ram[3539] = 8'h00;
    ff_ram[3540] = 8'h00;
    ff_ram[3541] = 8'h00;
    ff_ram[3542] = 8'h00;
    ff_ram[3543] = 8'h00;
    ff_ram[3544] = 8'h00;
    ff_ram[3545] = 8'h00;
    ff_ram[3546] = 8'h00;
    ff_ram[3547] = 8'h00;
    ff_ram[3548] = 8'h00;
    ff_ram[3549] = 8'h00;
    ff_ram[3550] = 8'h00;
    ff_ram[3551] = 8'h00;
    ff_ram[3552] = 8'h00;
    ff_ram[3553] = 8'h00;
    ff_ram[3554] = 8'h00;
    ff_ram[3555] = 8'h00;
    ff_ram[3556] = 8'h00;
    ff_ram[3557] = 8'h00;
    ff_ram[3558] = 8'h00;
    ff_ram[3559] = 8'h00;
    ff_ram[3560] = 8'h00;
    ff_ram[3561] = 8'h00;
    ff_ram[3562] = 8'h00;
    ff_ram[3563] = 8'h00;
    ff_ram[3564] = 8'h00;
    ff_ram[3565] = 8'h00;
    ff_ram[3566] = 8'h00;
    ff_ram[3567] = 8'h00;
    ff_ram[3568] = 8'h00;
    ff_ram[3569] = 8'h00;
    ff_ram[3570] = 8'h00;
    ff_ram[3571] = 8'h00;
    ff_ram[3572] = 8'h00;
    ff_ram[3573] = 8'h00;
    ff_ram[3574] = 8'h00;
    ff_ram[3575] = 8'h00;
    ff_ram[3576] = 8'h00;
    ff_ram[3577] = 8'h00;
    ff_ram[3578] = 8'h00;
    ff_ram[3579] = 8'h00;
    ff_ram[3580] = 8'h00;
    ff_ram[3581] = 8'h00;
    ff_ram[3582] = 8'h00;
    ff_ram[3583] = 8'h00;
    ff_ram[3584] = 8'h00;
    ff_ram[3585] = 8'h00;
    ff_ram[3586] = 8'h00;
    ff_ram[3587] = 8'h00;
    ff_ram[3588] = 8'h00;
    ff_ram[3589] = 8'h00;
    ff_ram[3590] = 8'h00;
    ff_ram[3591] = 8'h00;
    ff_ram[3592] = 8'h00;
    ff_ram[3593] = 8'h00;
    ff_ram[3594] = 8'h00;
    ff_ram[3595] = 8'h00;
    ff_ram[3596] = 8'h00;
    ff_ram[3597] = 8'h00;
    ff_ram[3598] = 8'h00;
    ff_ram[3599] = 8'h00;
    ff_ram[3600] = 8'h00;
    ff_ram[3601] = 8'h00;
    ff_ram[3602] = 8'h00;
    ff_ram[3603] = 8'h00;
    ff_ram[3604] = 8'h00;
    ff_ram[3605] = 8'h00;
    ff_ram[3606] = 8'h00;
    ff_ram[3607] = 8'h00;
    ff_ram[3608] = 8'h00;
    ff_ram[3609] = 8'h00;
    ff_ram[3610] = 8'h00;
    ff_ram[3611] = 8'h00;
    ff_ram[3612] = 8'h00;
    ff_ram[3613] = 8'h00;
    ff_ram[3614] = 8'h00;
    ff_ram[3615] = 8'h00;
    ff_ram[3616] = 8'h00;
    ff_ram[3617] = 8'h00;
    ff_ram[3618] = 8'h00;
    ff_ram[3619] = 8'h00;
    ff_ram[3620] = 8'h00;
    ff_ram[3621] = 8'h00;
    ff_ram[3622] = 8'h00;
    ff_ram[3623] = 8'h00;
    ff_ram[3624] = 8'h00;
    ff_ram[3625] = 8'h00;
    ff_ram[3626] = 8'h00;
    ff_ram[3627] = 8'h00;
    ff_ram[3628] = 8'h00;
    ff_ram[3629] = 8'h00;
    ff_ram[3630] = 8'h00;
    ff_ram[3631] = 8'h00;
    ff_ram[3632] = 8'h00;
    ff_ram[3633] = 8'h00;
    ff_ram[3634] = 8'h00;
    ff_ram[3635] = 8'h00;
    ff_ram[3636] = 8'h00;
    ff_ram[3637] = 8'h00;
    ff_ram[3638] = 8'h00;
    ff_ram[3639] = 8'h00;
    ff_ram[3640] = 8'h00;
    ff_ram[3641] = 8'h00;
    ff_ram[3642] = 8'h00;
    ff_ram[3643] = 8'h00;
    ff_ram[3644] = 8'h00;
    ff_ram[3645] = 8'h00;
    ff_ram[3646] = 8'h00;
    ff_ram[3647] = 8'h00;
    ff_ram[3648] = 8'h00;
    ff_ram[3649] = 8'h00;
    ff_ram[3650] = 8'h00;
    ff_ram[3651] = 8'h00;
    ff_ram[3652] = 8'h00;
    ff_ram[3653] = 8'h00;
    ff_ram[3654] = 8'h00;
    ff_ram[3655] = 8'h00;
    ff_ram[3656] = 8'h00;
    ff_ram[3657] = 8'h00;
    ff_ram[3658] = 8'h00;
    ff_ram[3659] = 8'h00;
    ff_ram[3660] = 8'h00;
    ff_ram[3661] = 8'h00;
    ff_ram[3662] = 8'h00;
    ff_ram[3663] = 8'h00;
    ff_ram[3664] = 8'h00;
    ff_ram[3665] = 8'h00;
    ff_ram[3666] = 8'h00;
    ff_ram[3667] = 8'h00;
    ff_ram[3668] = 8'h00;
    ff_ram[3669] = 8'h00;
    ff_ram[3670] = 8'h00;
    ff_ram[3671] = 8'h00;
    ff_ram[3672] = 8'h00;
    ff_ram[3673] = 8'h00;
    ff_ram[3674] = 8'h00;
    ff_ram[3675] = 8'h00;
    ff_ram[3676] = 8'h00;
    ff_ram[3677] = 8'h00;
    ff_ram[3678] = 8'h00;
    ff_ram[3679] = 8'h00;
    ff_ram[3680] = 8'h00;
    ff_ram[3681] = 8'h00;
    ff_ram[3682] = 8'h00;
    ff_ram[3683] = 8'h00;
    ff_ram[3684] = 8'h00;
    ff_ram[3685] = 8'h00;
    ff_ram[3686] = 8'h00;
    ff_ram[3687] = 8'h00;
    ff_ram[3688] = 8'h00;
    ff_ram[3689] = 8'h00;
    ff_ram[3690] = 8'h00;
    ff_ram[3691] = 8'h00;
    ff_ram[3692] = 8'h00;
    ff_ram[3693] = 8'h00;
    ff_ram[3694] = 8'h00;
    ff_ram[3695] = 8'h00;
    ff_ram[3696] = 8'h00;
    ff_ram[3697] = 8'h00;
    ff_ram[3698] = 8'h00;
    ff_ram[3699] = 8'h00;
    ff_ram[3700] = 8'h00;
    ff_ram[3701] = 8'h00;
    ff_ram[3702] = 8'h00;
    ff_ram[3703] = 8'h00;
    ff_ram[3704] = 8'h00;
    ff_ram[3705] = 8'h00;
    ff_ram[3706] = 8'h00;
    ff_ram[3707] = 8'h00;
    ff_ram[3708] = 8'h00;
    ff_ram[3709] = 8'h00;
    ff_ram[3710] = 8'h00;
    ff_ram[3711] = 8'h00;
    ff_ram[3712] = 8'h00;
    ff_ram[3713] = 8'h00;
    ff_ram[3714] = 8'h00;
    ff_ram[3715] = 8'h00;
    ff_ram[3716] = 8'h00;
    ff_ram[3717] = 8'h00;
    ff_ram[3718] = 8'h00;
    ff_ram[3719] = 8'h00;
    ff_ram[3720] = 8'h00;
    ff_ram[3721] = 8'h00;
    ff_ram[3722] = 8'h00;
    ff_ram[3723] = 8'h00;
    ff_ram[3724] = 8'h00;
    ff_ram[3725] = 8'h00;
    ff_ram[3726] = 8'h00;
    ff_ram[3727] = 8'h00;
    ff_ram[3728] = 8'h00;
    ff_ram[3729] = 8'h00;
    ff_ram[3730] = 8'h00;
    ff_ram[3731] = 8'h00;
    ff_ram[3732] = 8'h00;
    ff_ram[3733] = 8'h00;
    ff_ram[3734] = 8'h00;
    ff_ram[3735] = 8'h00;
    ff_ram[3736] = 8'h00;
    ff_ram[3737] = 8'h00;
    ff_ram[3738] = 8'h00;
    ff_ram[3739] = 8'h00;
    ff_ram[3740] = 8'h00;
    ff_ram[3741] = 8'h00;
    ff_ram[3742] = 8'h00;
    ff_ram[3743] = 8'h00;
    ff_ram[3744] = 8'h00;
    ff_ram[3745] = 8'h00;
    ff_ram[3746] = 8'h00;
    ff_ram[3747] = 8'h00;
    ff_ram[3748] = 8'h00;
    ff_ram[3749] = 8'h00;
    ff_ram[3750] = 8'h00;
    ff_ram[3751] = 8'h00;
    ff_ram[3752] = 8'h00;
    ff_ram[3753] = 8'h00;
    ff_ram[3754] = 8'h00;
    ff_ram[3755] = 8'h00;
    ff_ram[3756] = 8'h00;
    ff_ram[3757] = 8'h00;
    ff_ram[3758] = 8'h00;
    ff_ram[3759] = 8'h00;
    ff_ram[3760] = 8'h00;
    ff_ram[3761] = 8'h00;
    ff_ram[3762] = 8'h00;
    ff_ram[3763] = 8'h00;
    ff_ram[3764] = 8'h00;
    ff_ram[3765] = 8'h00;
    ff_ram[3766] = 8'h00;
    ff_ram[3767] = 8'h00;
    ff_ram[3768] = 8'h00;
    ff_ram[3769] = 8'h00;
    ff_ram[3770] = 8'h00;
    ff_ram[3771] = 8'h00;
    ff_ram[3772] = 8'h00;
    ff_ram[3773] = 8'h00;
    ff_ram[3774] = 8'h00;
    ff_ram[3775] = 8'h00;
    ff_ram[3776] = 8'h00;
    ff_ram[3777] = 8'h00;
    ff_ram[3778] = 8'h00;
    ff_ram[3779] = 8'h00;
    ff_ram[3780] = 8'h00;
    ff_ram[3781] = 8'h00;
    ff_ram[3782] = 8'h00;
    ff_ram[3783] = 8'h00;
    ff_ram[3784] = 8'h00;
    ff_ram[3785] = 8'h00;
    ff_ram[3786] = 8'h00;
    ff_ram[3787] = 8'h00;
    ff_ram[3788] = 8'h00;
    ff_ram[3789] = 8'h00;
    ff_ram[3790] = 8'h00;
    ff_ram[3791] = 8'h00;
    ff_ram[3792] = 8'h00;
    ff_ram[3793] = 8'h00;
    ff_ram[3794] = 8'h00;
    ff_ram[3795] = 8'h00;
    ff_ram[3796] = 8'h00;
    ff_ram[3797] = 8'h00;
    ff_ram[3798] = 8'h00;
    ff_ram[3799] = 8'h00;
    ff_ram[3800] = 8'h00;
    ff_ram[3801] = 8'h00;
    ff_ram[3802] = 8'h00;
    ff_ram[3803] = 8'h00;
    ff_ram[3804] = 8'h00;
    ff_ram[3805] = 8'h00;
    ff_ram[3806] = 8'h00;
    ff_ram[3807] = 8'h00;
    ff_ram[3808] = 8'h00;
    ff_ram[3809] = 8'h00;
    ff_ram[3810] = 8'h00;
    ff_ram[3811] = 8'h00;
    ff_ram[3812] = 8'h00;
    ff_ram[3813] = 8'h00;
    ff_ram[3814] = 8'h00;
    ff_ram[3815] = 8'h00;
    ff_ram[3816] = 8'h00;
    ff_ram[3817] = 8'h00;
    ff_ram[3818] = 8'h00;
    ff_ram[3819] = 8'h00;
    ff_ram[3820] = 8'h00;
    ff_ram[3821] = 8'h00;
    ff_ram[3822] = 8'h00;
    ff_ram[3823] = 8'h00;
    ff_ram[3824] = 8'h00;
    ff_ram[3825] = 8'h00;
    ff_ram[3826] = 8'h00;
    ff_ram[3827] = 8'h00;
    ff_ram[3828] = 8'h00;
    ff_ram[3829] = 8'h00;
    ff_ram[3830] = 8'h00;
    ff_ram[3831] = 8'h00;
    ff_ram[3832] = 8'h00;
    ff_ram[3833] = 8'h00;
    ff_ram[3834] = 8'h00;
    ff_ram[3835] = 8'h00;
    ff_ram[3836] = 8'h00;
    ff_ram[3837] = 8'h00;
    ff_ram[3838] = 8'h00;
    ff_ram[3839] = 8'h00;
    ff_ram[3840] = 8'h00;
    ff_ram[3841] = 8'h00;
    ff_ram[3842] = 8'h00;
    ff_ram[3843] = 8'h00;
    ff_ram[3844] = 8'h00;
    ff_ram[3845] = 8'h00;
    ff_ram[3846] = 8'h00;
    ff_ram[3847] = 8'h00;
    ff_ram[3848] = 8'h00;
    ff_ram[3849] = 8'h00;
    ff_ram[3850] = 8'h00;
    ff_ram[3851] = 8'h00;
    ff_ram[3852] = 8'h00;
    ff_ram[3853] = 8'h00;
    ff_ram[3854] = 8'h00;
    ff_ram[3855] = 8'h00;
    ff_ram[3856] = 8'h00;
    ff_ram[3857] = 8'h00;
    ff_ram[3858] = 8'h00;
    ff_ram[3859] = 8'h00;
    ff_ram[3860] = 8'h00;
    ff_ram[3861] = 8'h00;
    ff_ram[3862] = 8'h00;
    ff_ram[3863] = 8'h00;
    ff_ram[3864] = 8'h00;
    ff_ram[3865] = 8'h00;
    ff_ram[3866] = 8'h00;
    ff_ram[3867] = 8'h00;
    ff_ram[3868] = 8'h00;
    ff_ram[3869] = 8'h00;
    ff_ram[3870] = 8'h00;
    ff_ram[3871] = 8'h00;
    ff_ram[3872] = 8'h00;
    ff_ram[3873] = 8'h00;
    ff_ram[3874] = 8'h00;
    ff_ram[3875] = 8'h00;
    ff_ram[3876] = 8'h00;
    ff_ram[3877] = 8'h00;
    ff_ram[3878] = 8'h00;
    ff_ram[3879] = 8'h00;
    ff_ram[3880] = 8'h00;
    ff_ram[3881] = 8'h00;
    ff_ram[3882] = 8'h00;
    ff_ram[3883] = 8'h00;
    ff_ram[3884] = 8'h00;
    ff_ram[3885] = 8'h00;
    ff_ram[3886] = 8'h00;
    ff_ram[3887] = 8'h00;
    ff_ram[3888] = 8'h00;
    ff_ram[3889] = 8'h00;
    ff_ram[3890] = 8'h00;
    ff_ram[3891] = 8'h00;
    ff_ram[3892] = 8'h00;
    ff_ram[3893] = 8'h00;
    ff_ram[3894] = 8'h00;
    ff_ram[3895] = 8'h00;
    ff_ram[3896] = 8'h00;
    ff_ram[3897] = 8'h00;
    ff_ram[3898] = 8'h00;
    ff_ram[3899] = 8'h00;
    ff_ram[3900] = 8'h00;
    ff_ram[3901] = 8'h00;
    ff_ram[3902] = 8'h00;
    ff_ram[3903] = 8'h00;
    ff_ram[3904] = 8'h00;
    ff_ram[3905] = 8'h00;
    ff_ram[3906] = 8'h00;
    ff_ram[3907] = 8'h00;
    ff_ram[3908] = 8'h00;
    ff_ram[3909] = 8'h00;
    ff_ram[3910] = 8'h00;
    ff_ram[3911] = 8'h00;
    ff_ram[3912] = 8'h00;
    ff_ram[3913] = 8'h00;
    ff_ram[3914] = 8'h00;
    ff_ram[3915] = 8'h00;
    ff_ram[3916] = 8'h00;
    ff_ram[3917] = 8'h00;
    ff_ram[3918] = 8'h00;
    ff_ram[3919] = 8'h00;
    ff_ram[3920] = 8'h00;
    ff_ram[3921] = 8'h00;
    ff_ram[3922] = 8'h00;
    ff_ram[3923] = 8'h00;
    ff_ram[3924] = 8'h00;
    ff_ram[3925] = 8'h00;
    ff_ram[3926] = 8'h00;
    ff_ram[3927] = 8'h00;
    ff_ram[3928] = 8'h00;
    ff_ram[3929] = 8'h00;
    ff_ram[3930] = 8'h00;
    ff_ram[3931] = 8'h00;
    ff_ram[3932] = 8'h00;
    ff_ram[3933] = 8'h00;
    ff_ram[3934] = 8'h00;
    ff_ram[3935] = 8'h00;
    ff_ram[3936] = 8'h00;
    ff_ram[3937] = 8'h00;
    ff_ram[3938] = 8'h00;
    ff_ram[3939] = 8'h00;
    ff_ram[3940] = 8'h00;
    ff_ram[3941] = 8'h00;
    ff_ram[3942] = 8'h00;
    ff_ram[3943] = 8'h00;
    ff_ram[3944] = 8'h00;
    ff_ram[3945] = 8'h00;
    ff_ram[3946] = 8'h00;
    ff_ram[3947] = 8'h00;
    ff_ram[3948] = 8'h00;
    ff_ram[3949] = 8'h00;
    ff_ram[3950] = 8'h00;
    ff_ram[3951] = 8'h00;
    ff_ram[3952] = 8'h00;
    ff_ram[3953] = 8'h00;
    ff_ram[3954] = 8'h00;
    ff_ram[3955] = 8'h00;
    ff_ram[3956] = 8'h00;
    ff_ram[3957] = 8'h00;
    ff_ram[3958] = 8'h00;
    ff_ram[3959] = 8'h00;
    ff_ram[3960] = 8'h00;
    ff_ram[3961] = 8'h00;
    ff_ram[3962] = 8'h00;
    ff_ram[3963] = 8'h00;
    ff_ram[3964] = 8'h00;
    ff_ram[3965] = 8'h00;
    ff_ram[3966] = 8'h00;
    ff_ram[3967] = 8'h00;
    ff_ram[3968] = 8'h00;
    ff_ram[3969] = 8'h00;
    ff_ram[3970] = 8'h00;
    ff_ram[3971] = 8'h00;
    ff_ram[3972] = 8'h00;
    ff_ram[3973] = 8'h00;
    ff_ram[3974] = 8'h00;
    ff_ram[3975] = 8'h00;
    ff_ram[3976] = 8'h00;
    ff_ram[3977] = 8'h00;
    ff_ram[3978] = 8'h00;
    ff_ram[3979] = 8'h00;
    ff_ram[3980] = 8'h00;
    ff_ram[3981] = 8'h00;
    ff_ram[3982] = 8'h00;
    ff_ram[3983] = 8'h00;
    ff_ram[3984] = 8'h00;
    ff_ram[3985] = 8'h00;
    ff_ram[3986] = 8'h00;
    ff_ram[3987] = 8'h00;
    ff_ram[3988] = 8'h00;
    ff_ram[3989] = 8'h00;
    ff_ram[3990] = 8'h00;
    ff_ram[3991] = 8'h00;
    ff_ram[3992] = 8'h00;
    ff_ram[3993] = 8'h00;
    ff_ram[3994] = 8'h00;
    ff_ram[3995] = 8'h00;
    ff_ram[3996] = 8'h00;
    ff_ram[3997] = 8'h00;
    ff_ram[3998] = 8'h00;
    ff_ram[3999] = 8'h00;
    ff_ram[4000] = 8'h00;
    ff_ram[4001] = 8'h00;
    ff_ram[4002] = 8'h00;
    ff_ram[4003] = 8'h00;
    ff_ram[4004] = 8'h00;
    ff_ram[4005] = 8'h00;
    ff_ram[4006] = 8'h00;
    ff_ram[4007] = 8'h00;
    ff_ram[4008] = 8'h00;
    ff_ram[4009] = 8'h00;
    ff_ram[4010] = 8'h00;
    ff_ram[4011] = 8'h00;
    ff_ram[4012] = 8'h00;
    ff_ram[4013] = 8'h00;
    ff_ram[4014] = 8'h00;
    ff_ram[4015] = 8'h00;
    ff_ram[4016] = 8'h00;
    ff_ram[4017] = 8'h00;
    ff_ram[4018] = 8'h00;
    ff_ram[4019] = 8'h00;
    ff_ram[4020] = 8'h00;
    ff_ram[4021] = 8'h00;
    ff_ram[4022] = 8'h00;
    ff_ram[4023] = 8'h00;
    ff_ram[4024] = 8'h00;
    ff_ram[4025] = 8'h00;
    ff_ram[4026] = 8'h00;
    ff_ram[4027] = 8'h00;
    ff_ram[4028] = 8'h00;
    ff_ram[4029] = 8'h00;
    ff_ram[4030] = 8'h00;
    ff_ram[4031] = 8'h00;
    ff_ram[4032] = 8'h00;
    ff_ram[4033] = 8'h00;
    ff_ram[4034] = 8'h00;
    ff_ram[4035] = 8'h00;
    ff_ram[4036] = 8'h00;
    ff_ram[4037] = 8'h00;
    ff_ram[4038] = 8'h00;
    ff_ram[4039] = 8'h00;
    ff_ram[4040] = 8'h00;
    ff_ram[4041] = 8'h00;
    ff_ram[4042] = 8'h00;
    ff_ram[4043] = 8'h00;
    ff_ram[4044] = 8'h00;
    ff_ram[4045] = 8'h00;
    ff_ram[4046] = 8'h00;
    ff_ram[4047] = 8'h00;
    ff_ram[4048] = 8'h00;
    ff_ram[4049] = 8'h00;
    ff_ram[4050] = 8'h00;
    ff_ram[4051] = 8'h00;
    ff_ram[4052] = 8'h00;
    ff_ram[4053] = 8'h00;
    ff_ram[4054] = 8'h00;
    ff_ram[4055] = 8'h00;
    ff_ram[4056] = 8'h00;
    ff_ram[4057] = 8'h00;
    ff_ram[4058] = 8'h00;
    ff_ram[4059] = 8'h00;
    ff_ram[4060] = 8'h00;
    ff_ram[4061] = 8'h00;
    ff_ram[4062] = 8'h00;
    ff_ram[4063] = 8'h00;
    ff_ram[4064] = 8'h00;
    ff_ram[4065] = 8'h00;
    ff_ram[4066] = 8'h00;
    ff_ram[4067] = 8'h00;
    ff_ram[4068] = 8'h00;
    ff_ram[4069] = 8'h00;
    ff_ram[4070] = 8'h00;
    ff_ram[4071] = 8'h00;
    ff_ram[4072] = 8'h00;
    ff_ram[4073] = 8'h00;
    ff_ram[4074] = 8'h00;
    ff_ram[4075] = 8'h00;
    ff_ram[4076] = 8'h00;
    ff_ram[4077] = 8'h00;
    ff_ram[4078] = 8'h00;
    ff_ram[4079] = 8'h00;
    ff_ram[4080] = 8'h00;
    ff_ram[4081] = 8'h00;
    ff_ram[4082] = 8'h00;
    ff_ram[4083] = 8'h00;
    ff_ram[4084] = 8'h00;
    ff_ram[4085] = 8'h00;
    ff_ram[4086] = 8'h00;
    ff_ram[4087] = 8'h00;
    ff_ram[4088] = 8'h00;
    ff_ram[4089] = 8'h00;
    ff_ram[4090] = 8'h00;
    ff_ram[4091] = 8'h00;
    ff_ram[4092] = 8'h00;
    ff_ram[4093] = 8'h00;
    ff_ram[4094] = 8'h00;
    ff_ram[4095] = 8'h00;
    ff_ram[4096] = 8'h00;
    ff_ram[4097] = 8'h00;
    ff_ram[4098] = 8'h00;
    ff_ram[4099] = 8'h00;
    ff_ram[4100] = 8'h00;
    ff_ram[4101] = 8'h00;
    ff_ram[4102] = 8'h00;
    ff_ram[4103] = 8'h00;
    ff_ram[4104] = 8'h00;
    ff_ram[4105] = 8'h00;
    ff_ram[4106] = 8'h00;
    ff_ram[4107] = 8'h00;
    ff_ram[4108] = 8'h00;
    ff_ram[4109] = 8'h00;
    ff_ram[4110] = 8'h00;
    ff_ram[4111] = 8'h00;
    ff_ram[4112] = 8'h00;
    ff_ram[4113] = 8'h00;
    ff_ram[4114] = 8'h00;
    ff_ram[4115] = 8'h00;
    ff_ram[4116] = 8'h00;
    ff_ram[4117] = 8'h00;
    ff_ram[4118] = 8'h00;
    ff_ram[4119] = 8'h00;
    ff_ram[4120] = 8'h00;
    ff_ram[4121] = 8'h00;
    ff_ram[4122] = 8'h00;
    ff_ram[4123] = 8'h00;
    ff_ram[4124] = 8'h00;
    ff_ram[4125] = 8'h00;
    ff_ram[4126] = 8'h00;
    ff_ram[4127] = 8'h00;
    ff_ram[4128] = 8'h00;
    ff_ram[4129] = 8'h00;
    ff_ram[4130] = 8'h00;
    ff_ram[4131] = 8'h00;
    ff_ram[4132] = 8'h00;
    ff_ram[4133] = 8'h00;
    ff_ram[4134] = 8'h00;
    ff_ram[4135] = 8'h00;
    ff_ram[4136] = 8'h00;
    ff_ram[4137] = 8'h00;
    ff_ram[4138] = 8'h00;
    ff_ram[4139] = 8'h00;
    ff_ram[4140] = 8'h00;
    ff_ram[4141] = 8'h00;
    ff_ram[4142] = 8'h00;
    ff_ram[4143] = 8'h00;
    ff_ram[4144] = 8'h00;
    ff_ram[4145] = 8'h00;
    ff_ram[4146] = 8'h00;
    ff_ram[4147] = 8'h00;
    ff_ram[4148] = 8'h00;
    ff_ram[4149] = 8'h00;
    ff_ram[4150] = 8'h00;
    ff_ram[4151] = 8'h00;
    ff_ram[4152] = 8'h00;
    ff_ram[4153] = 8'h00;
    ff_ram[4154] = 8'h00;
    ff_ram[4155] = 8'h00;
    ff_ram[4156] = 8'h00;
    ff_ram[4157] = 8'h00;
    ff_ram[4158] = 8'h00;
    ff_ram[4159] = 8'h00;
    ff_ram[4160] = 8'h00;
    ff_ram[4161] = 8'h00;
    ff_ram[4162] = 8'h00;
    ff_ram[4163] = 8'h00;
    ff_ram[4164] = 8'h00;
    ff_ram[4165] = 8'h00;
    ff_ram[4166] = 8'h00;
    ff_ram[4167] = 8'h00;
    ff_ram[4168] = 8'h00;
    ff_ram[4169] = 8'h00;
    ff_ram[4170] = 8'h00;
    ff_ram[4171] = 8'h00;
    ff_ram[4172] = 8'h00;
    ff_ram[4173] = 8'h00;
    ff_ram[4174] = 8'h00;
    ff_ram[4175] = 8'h00;
    ff_ram[4176] = 8'h00;
    ff_ram[4177] = 8'h00;
    ff_ram[4178] = 8'h00;
    ff_ram[4179] = 8'h00;
    ff_ram[4180] = 8'h00;
    ff_ram[4181] = 8'h00;
    ff_ram[4182] = 8'h00;
    ff_ram[4183] = 8'h00;
    ff_ram[4184] = 8'h00;
    ff_ram[4185] = 8'h00;
    ff_ram[4186] = 8'h00;
    ff_ram[4187] = 8'h00;
    ff_ram[4188] = 8'h00;
    ff_ram[4189] = 8'h00;
    ff_ram[4190] = 8'h00;
    ff_ram[4191] = 8'h00;
    ff_ram[4192] = 8'h00;
    ff_ram[4193] = 8'h00;
    ff_ram[4194] = 8'h00;
    ff_ram[4195] = 8'h00;
    ff_ram[4196] = 8'h00;
    ff_ram[4197] = 8'h00;
    ff_ram[4198] = 8'h00;
    ff_ram[4199] = 8'h00;
    ff_ram[4200] = 8'h00;
    ff_ram[4201] = 8'h00;
    ff_ram[4202] = 8'h00;
    ff_ram[4203] = 8'h00;
    ff_ram[4204] = 8'h00;
    ff_ram[4205] = 8'h00;
    ff_ram[4206] = 8'h00;
    ff_ram[4207] = 8'h00;
    ff_ram[4208] = 8'h00;
    ff_ram[4209] = 8'h00;
    ff_ram[4210] = 8'h00;
    ff_ram[4211] = 8'h00;
    ff_ram[4212] = 8'h00;
    ff_ram[4213] = 8'h00;
    ff_ram[4214] = 8'h00;
    ff_ram[4215] = 8'h00;
    ff_ram[4216] = 8'h00;
    ff_ram[4217] = 8'h00;
    ff_ram[4218] = 8'h00;
    ff_ram[4219] = 8'h00;
    ff_ram[4220] = 8'h00;
    ff_ram[4221] = 8'h00;
    ff_ram[4222] = 8'h00;
    ff_ram[4223] = 8'h00;
    ff_ram[4224] = 8'h00;
    ff_ram[4225] = 8'h00;
    ff_ram[4226] = 8'h00;
    ff_ram[4227] = 8'h00;
    ff_ram[4228] = 8'h00;
    ff_ram[4229] = 8'h00;
    ff_ram[4230] = 8'h00;
    ff_ram[4231] = 8'h00;
    ff_ram[4232] = 8'h00;
    ff_ram[4233] = 8'h00;
    ff_ram[4234] = 8'h00;
    ff_ram[4235] = 8'h00;
    ff_ram[4236] = 8'h00;
    ff_ram[4237] = 8'h00;
    ff_ram[4238] = 8'h00;
    ff_ram[4239] = 8'h00;
    ff_ram[4240] = 8'h00;
    ff_ram[4241] = 8'h00;
    ff_ram[4242] = 8'h00;
    ff_ram[4243] = 8'h00;
    ff_ram[4244] = 8'h00;
    ff_ram[4245] = 8'h00;
    ff_ram[4246] = 8'h00;
    ff_ram[4247] = 8'h00;
    ff_ram[4248] = 8'h00;
    ff_ram[4249] = 8'h00;
    ff_ram[4250] = 8'h00;
    ff_ram[4251] = 8'h00;
    ff_ram[4252] = 8'h00;
    ff_ram[4253] = 8'h00;
    ff_ram[4254] = 8'h00;
    ff_ram[4255] = 8'h00;
    ff_ram[4256] = 8'h00;
    ff_ram[4257] = 8'h00;
    ff_ram[4258] = 8'h00;
    ff_ram[4259] = 8'h00;
    ff_ram[4260] = 8'h00;
    ff_ram[4261] = 8'h00;
    ff_ram[4262] = 8'h00;
    ff_ram[4263] = 8'h00;
    ff_ram[4264] = 8'h00;
    ff_ram[4265] = 8'h00;
    ff_ram[4266] = 8'h00;
    ff_ram[4267] = 8'h00;
    ff_ram[4268] = 8'h00;
    ff_ram[4269] = 8'h00;
    ff_ram[4270] = 8'h00;
    ff_ram[4271] = 8'h00;
    ff_ram[4272] = 8'h00;
    ff_ram[4273] = 8'h00;
    ff_ram[4274] = 8'h00;
    ff_ram[4275] = 8'h00;
    ff_ram[4276] = 8'h00;
    ff_ram[4277] = 8'h00;
    ff_ram[4278] = 8'h00;
    ff_ram[4279] = 8'h00;
    ff_ram[4280] = 8'h00;
    ff_ram[4281] = 8'h00;
    ff_ram[4282] = 8'h00;
    ff_ram[4283] = 8'h00;
    ff_ram[4284] = 8'h00;
    ff_ram[4285] = 8'h00;
    ff_ram[4286] = 8'h00;
    ff_ram[4287] = 8'h00;
    ff_ram[4288] = 8'h00;
    ff_ram[4289] = 8'h00;
    ff_ram[4290] = 8'h00;
    ff_ram[4291] = 8'h00;
    ff_ram[4292] = 8'h00;
    ff_ram[4293] = 8'h00;
    ff_ram[4294] = 8'h00;
    ff_ram[4295] = 8'h00;
    ff_ram[4296] = 8'h00;
    ff_ram[4297] = 8'h00;
    ff_ram[4298] = 8'h00;
    ff_ram[4299] = 8'h00;
    ff_ram[4300] = 8'h00;
    ff_ram[4301] = 8'h00;
    ff_ram[4302] = 8'h00;
    ff_ram[4303] = 8'h00;
    ff_ram[4304] = 8'h00;
    ff_ram[4305] = 8'h00;
    ff_ram[4306] = 8'h00;
    ff_ram[4307] = 8'h00;
    ff_ram[4308] = 8'h00;
    ff_ram[4309] = 8'h00;
    ff_ram[4310] = 8'h00;
    ff_ram[4311] = 8'h00;
    ff_ram[4312] = 8'h00;
    ff_ram[4313] = 8'h00;
    ff_ram[4314] = 8'h00;
    ff_ram[4315] = 8'h00;
    ff_ram[4316] = 8'h00;
    ff_ram[4317] = 8'h00;
    ff_ram[4318] = 8'h00;
    ff_ram[4319] = 8'h00;
    ff_ram[4320] = 8'h00;
    ff_ram[4321] = 8'h00;
    ff_ram[4322] = 8'h00;
    ff_ram[4323] = 8'h00;
    ff_ram[4324] = 8'h00;
    ff_ram[4325] = 8'h00;
    ff_ram[4326] = 8'h00;
    ff_ram[4327] = 8'h00;
    ff_ram[4328] = 8'h00;
    ff_ram[4329] = 8'h00;
    ff_ram[4330] = 8'h00;
    ff_ram[4331] = 8'h00;
    ff_ram[4332] = 8'h00;
    ff_ram[4333] = 8'h00;
    ff_ram[4334] = 8'h00;
    ff_ram[4335] = 8'h00;
    ff_ram[4336] = 8'h00;
    ff_ram[4337] = 8'h00;
    ff_ram[4338] = 8'h00;
    ff_ram[4339] = 8'h00;
    ff_ram[4340] = 8'h00;
    ff_ram[4341] = 8'h00;
    ff_ram[4342] = 8'h00;
    ff_ram[4343] = 8'h00;
    ff_ram[4344] = 8'h00;
    ff_ram[4345] = 8'h00;
    ff_ram[4346] = 8'h00;
    ff_ram[4347] = 8'h00;
    ff_ram[4348] = 8'h00;
    ff_ram[4349] = 8'h00;
    ff_ram[4350] = 8'h00;
    ff_ram[4351] = 8'h00;
    ff_ram[4352] = 8'h00;
    ff_ram[4353] = 8'h00;
    ff_ram[4354] = 8'h00;
    ff_ram[4355] = 8'h00;
    ff_ram[4356] = 8'h00;
    ff_ram[4357] = 8'h00;
    ff_ram[4358] = 8'h00;
    ff_ram[4359] = 8'h00;
    ff_ram[4360] = 8'h00;
    ff_ram[4361] = 8'h00;
    ff_ram[4362] = 8'h00;
    ff_ram[4363] = 8'h00;
    ff_ram[4364] = 8'h00;
    ff_ram[4365] = 8'h00;
    ff_ram[4366] = 8'h00;
    ff_ram[4367] = 8'h00;
    ff_ram[4368] = 8'h00;
    ff_ram[4369] = 8'h00;
    ff_ram[4370] = 8'h00;
    ff_ram[4371] = 8'h00;
    ff_ram[4372] = 8'h00;
    ff_ram[4373] = 8'h00;
    ff_ram[4374] = 8'h00;
    ff_ram[4375] = 8'h00;
    ff_ram[4376] = 8'h00;
    ff_ram[4377] = 8'h00;
    ff_ram[4378] = 8'h00;
    ff_ram[4379] = 8'h00;
    ff_ram[4380] = 8'h00;
    ff_ram[4381] = 8'h00;
    ff_ram[4382] = 8'h00;
    ff_ram[4383] = 8'h00;
    ff_ram[4384] = 8'h00;
    ff_ram[4385] = 8'h00;
    ff_ram[4386] = 8'h00;
    ff_ram[4387] = 8'h00;
    ff_ram[4388] = 8'h00;
    ff_ram[4389] = 8'h00;
    ff_ram[4390] = 8'h00;
    ff_ram[4391] = 8'h00;
    ff_ram[4392] = 8'h00;
    ff_ram[4393] = 8'h00;
    ff_ram[4394] = 8'h00;
    ff_ram[4395] = 8'h00;
    ff_ram[4396] = 8'h00;
    ff_ram[4397] = 8'h00;
    ff_ram[4398] = 8'h00;
    ff_ram[4399] = 8'h00;
    ff_ram[4400] = 8'h00;
    ff_ram[4401] = 8'h00;
    ff_ram[4402] = 8'h00;
    ff_ram[4403] = 8'h00;
    ff_ram[4404] = 8'h00;
    ff_ram[4405] = 8'h00;
    ff_ram[4406] = 8'h00;
    ff_ram[4407] = 8'h00;
    ff_ram[4408] = 8'h00;
    ff_ram[4409] = 8'h00;
    ff_ram[4410] = 8'h00;
    ff_ram[4411] = 8'h00;
    ff_ram[4412] = 8'h00;
    ff_ram[4413] = 8'h00;
    ff_ram[4414] = 8'h00;
    ff_ram[4415] = 8'h00;
    ff_ram[4416] = 8'h00;
    ff_ram[4417] = 8'h00;
    ff_ram[4418] = 8'h00;
    ff_ram[4419] = 8'h00;
    ff_ram[4420] = 8'h00;
    ff_ram[4421] = 8'h00;
    ff_ram[4422] = 8'h00;
    ff_ram[4423] = 8'h00;
    ff_ram[4424] = 8'h00;
    ff_ram[4425] = 8'h00;
    ff_ram[4426] = 8'h00;
    ff_ram[4427] = 8'h00;
    ff_ram[4428] = 8'h00;
    ff_ram[4429] = 8'h00;
    ff_ram[4430] = 8'h00;
    ff_ram[4431] = 8'h00;
    ff_ram[4432] = 8'h00;
    ff_ram[4433] = 8'h00;
    ff_ram[4434] = 8'h00;
    ff_ram[4435] = 8'h00;
    ff_ram[4436] = 8'h00;
    ff_ram[4437] = 8'h00;
    ff_ram[4438] = 8'h00;
    ff_ram[4439] = 8'h00;
    ff_ram[4440] = 8'h00;
    ff_ram[4441] = 8'h00;
    ff_ram[4442] = 8'h00;
    ff_ram[4443] = 8'h00;
    ff_ram[4444] = 8'h00;
    ff_ram[4445] = 8'h00;
    ff_ram[4446] = 8'h00;
    ff_ram[4447] = 8'h00;
    ff_ram[4448] = 8'h00;
    ff_ram[4449] = 8'h00;
    ff_ram[4450] = 8'h00;
    ff_ram[4451] = 8'h00;
    ff_ram[4452] = 8'h00;
    ff_ram[4453] = 8'h00;
    ff_ram[4454] = 8'h00;
    ff_ram[4455] = 8'h00;
    ff_ram[4456] = 8'h00;
    ff_ram[4457] = 8'h00;
    ff_ram[4458] = 8'h00;
    ff_ram[4459] = 8'h00;
    ff_ram[4460] = 8'h00;
    ff_ram[4461] = 8'h00;
    ff_ram[4462] = 8'h00;
    ff_ram[4463] = 8'h00;
    ff_ram[4464] = 8'h00;
    ff_ram[4465] = 8'h00;
    ff_ram[4466] = 8'h00;
    ff_ram[4467] = 8'h00;
    ff_ram[4468] = 8'h00;
    ff_ram[4469] = 8'h00;
    ff_ram[4470] = 8'h00;
    ff_ram[4471] = 8'h00;
    ff_ram[4472] = 8'h00;
    ff_ram[4473] = 8'h00;
    ff_ram[4474] = 8'h00;
    ff_ram[4475] = 8'h00;
    ff_ram[4476] = 8'h00;
    ff_ram[4477] = 8'h00;
    ff_ram[4478] = 8'h00;
    ff_ram[4479] = 8'h00;
    ff_ram[4480] = 8'h00;
    ff_ram[4481] = 8'h00;
    ff_ram[4482] = 8'h00;
    ff_ram[4483] = 8'h00;
    ff_ram[4484] = 8'h00;
    ff_ram[4485] = 8'h00;
    ff_ram[4486] = 8'h00;
    ff_ram[4487] = 8'h00;
    ff_ram[4488] = 8'h00;
    ff_ram[4489] = 8'h00;
    ff_ram[4490] = 8'h00;
    ff_ram[4491] = 8'h00;
    ff_ram[4492] = 8'h00;
    ff_ram[4493] = 8'h00;
    ff_ram[4494] = 8'h00;
    ff_ram[4495] = 8'h00;
    ff_ram[4496] = 8'h00;
    ff_ram[4497] = 8'h00;
    ff_ram[4498] = 8'h00;
    ff_ram[4499] = 8'h00;
    ff_ram[4500] = 8'h00;
    ff_ram[4501] = 8'h00;
    ff_ram[4502] = 8'h00;
    ff_ram[4503] = 8'h00;
    ff_ram[4504] = 8'h00;
    ff_ram[4505] = 8'h00;
    ff_ram[4506] = 8'h00;
    ff_ram[4507] = 8'h00;
    ff_ram[4508] = 8'h00;
    ff_ram[4509] = 8'h00;
    ff_ram[4510] = 8'h00;
    ff_ram[4511] = 8'h00;
    ff_ram[4512] = 8'h00;
    ff_ram[4513] = 8'h00;
    ff_ram[4514] = 8'h00;
    ff_ram[4515] = 8'h00;
    ff_ram[4516] = 8'h00;
    ff_ram[4517] = 8'h00;
    ff_ram[4518] = 8'h00;
    ff_ram[4519] = 8'h00;
    ff_ram[4520] = 8'h00;
    ff_ram[4521] = 8'h00;
    ff_ram[4522] = 8'h00;
    ff_ram[4523] = 8'h00;
    ff_ram[4524] = 8'h00;
    ff_ram[4525] = 8'h00;
    ff_ram[4526] = 8'h00;
    ff_ram[4527] = 8'h00;
    ff_ram[4528] = 8'h00;
    ff_ram[4529] = 8'h00;
    ff_ram[4530] = 8'h00;
    ff_ram[4531] = 8'h00;
    ff_ram[4532] = 8'h00;
    ff_ram[4533] = 8'h00;
    ff_ram[4534] = 8'h00;
    ff_ram[4535] = 8'h00;
    ff_ram[4536] = 8'h00;
    ff_ram[4537] = 8'h00;
    ff_ram[4538] = 8'h00;
    ff_ram[4539] = 8'h00;
    ff_ram[4540] = 8'h00;
    ff_ram[4541] = 8'h00;
    ff_ram[4542] = 8'h00;
    ff_ram[4543] = 8'h00;
    ff_ram[4544] = 8'h00;
    ff_ram[4545] = 8'h00;
    ff_ram[4546] = 8'h00;
    ff_ram[4547] = 8'h00;
    ff_ram[4548] = 8'h00;
    ff_ram[4549] = 8'h00;
    ff_ram[4550] = 8'h00;
    ff_ram[4551] = 8'h00;
    ff_ram[4552] = 8'h00;
    ff_ram[4553] = 8'h00;
    ff_ram[4554] = 8'h00;
    ff_ram[4555] = 8'h00;
    ff_ram[4556] = 8'h00;
    ff_ram[4557] = 8'h00;
    ff_ram[4558] = 8'h00;
    ff_ram[4559] = 8'h00;
    ff_ram[4560] = 8'h00;
    ff_ram[4561] = 8'h00;
    ff_ram[4562] = 8'h00;
    ff_ram[4563] = 8'h00;
    ff_ram[4564] = 8'h00;
    ff_ram[4565] = 8'h00;
    ff_ram[4566] = 8'h00;
    ff_ram[4567] = 8'h00;
    ff_ram[4568] = 8'h00;
    ff_ram[4569] = 8'h00;
    ff_ram[4570] = 8'h00;
    ff_ram[4571] = 8'h00;
    ff_ram[4572] = 8'h00;
    ff_ram[4573] = 8'h00;
    ff_ram[4574] = 8'h00;
    ff_ram[4575] = 8'h00;
    ff_ram[4576] = 8'h00;
    ff_ram[4577] = 8'h00;
    ff_ram[4578] = 8'h00;
    ff_ram[4579] = 8'h00;
    ff_ram[4580] = 8'h00;
    ff_ram[4581] = 8'h00;
    ff_ram[4582] = 8'h00;
    ff_ram[4583] = 8'h00;
    ff_ram[4584] = 8'h00;
    ff_ram[4585] = 8'h00;
    ff_ram[4586] = 8'h00;
    ff_ram[4587] = 8'h00;
    ff_ram[4588] = 8'h00;
    ff_ram[4589] = 8'h00;
    ff_ram[4590] = 8'h00;
    ff_ram[4591] = 8'h00;
    ff_ram[4592] = 8'h00;
    ff_ram[4593] = 8'h00;
    ff_ram[4594] = 8'h00;
    ff_ram[4595] = 8'h00;
    ff_ram[4596] = 8'h00;
    ff_ram[4597] = 8'h00;
    ff_ram[4598] = 8'h00;
    ff_ram[4599] = 8'h00;
    ff_ram[4600] = 8'h00;
    ff_ram[4601] = 8'h00;
    ff_ram[4602] = 8'h00;
    ff_ram[4603] = 8'h00;
    ff_ram[4604] = 8'h00;
    ff_ram[4605] = 8'h00;
    ff_ram[4606] = 8'h00;
    ff_ram[4607] = 8'h00;
    ff_ram[4608] = 8'h00;
    ff_ram[4609] = 8'h00;
    ff_ram[4610] = 8'h00;
    ff_ram[4611] = 8'h00;
    ff_ram[4612] = 8'h00;
    ff_ram[4613] = 8'h00;
    ff_ram[4614] = 8'h00;
    ff_ram[4615] = 8'h00;
    ff_ram[4616] = 8'h00;
    ff_ram[4617] = 8'h00;
    ff_ram[4618] = 8'h00;
    ff_ram[4619] = 8'h00;
    ff_ram[4620] = 8'h00;
    ff_ram[4621] = 8'h00;
    ff_ram[4622] = 8'h00;
    ff_ram[4623] = 8'h00;
    ff_ram[4624] = 8'h00;
    ff_ram[4625] = 8'h00;
    ff_ram[4626] = 8'h00;
    ff_ram[4627] = 8'h00;
    ff_ram[4628] = 8'h00;
    ff_ram[4629] = 8'h00;
    ff_ram[4630] = 8'h00;
    ff_ram[4631] = 8'h00;
    ff_ram[4632] = 8'h00;
    ff_ram[4633] = 8'h00;
    ff_ram[4634] = 8'h00;
    ff_ram[4635] = 8'h00;
    ff_ram[4636] = 8'h00;
    ff_ram[4637] = 8'h00;
    ff_ram[4638] = 8'h00;
    ff_ram[4639] = 8'h00;
    ff_ram[4640] = 8'h00;
    ff_ram[4641] = 8'h00;
    ff_ram[4642] = 8'h00;
    ff_ram[4643] = 8'h00;
    ff_ram[4644] = 8'h00;
    ff_ram[4645] = 8'h00;
    ff_ram[4646] = 8'h00;
    ff_ram[4647] = 8'h00;
    ff_ram[4648] = 8'h00;
    ff_ram[4649] = 8'h00;
    ff_ram[4650] = 8'h00;
    ff_ram[4651] = 8'h00;
    ff_ram[4652] = 8'h00;
    ff_ram[4653] = 8'h00;
    ff_ram[4654] = 8'h00;
    ff_ram[4655] = 8'h00;
    ff_ram[4656] = 8'h00;
    ff_ram[4657] = 8'h00;
    ff_ram[4658] = 8'h00;
    ff_ram[4659] = 8'h00;
    ff_ram[4660] = 8'h00;
    ff_ram[4661] = 8'h00;
    ff_ram[4662] = 8'h00;
    ff_ram[4663] = 8'h00;
    ff_ram[4664] = 8'h00;
    ff_ram[4665] = 8'h00;
    ff_ram[4666] = 8'h00;
    ff_ram[4667] = 8'h00;
    ff_ram[4668] = 8'h00;
    ff_ram[4669] = 8'h00;
    ff_ram[4670] = 8'h00;
    ff_ram[4671] = 8'h00;
    ff_ram[4672] = 8'h00;
    ff_ram[4673] = 8'h00;
    ff_ram[4674] = 8'h00;
    ff_ram[4675] = 8'h00;
    ff_ram[4676] = 8'h00;
    ff_ram[4677] = 8'h00;
    ff_ram[4678] = 8'h00;
    ff_ram[4679] = 8'h00;
    ff_ram[4680] = 8'h00;
    ff_ram[4681] = 8'h00;
    ff_ram[4682] = 8'h00;
    ff_ram[4683] = 8'h00;
    ff_ram[4684] = 8'h00;
    ff_ram[4685] = 8'h00;
    ff_ram[4686] = 8'h00;
    ff_ram[4687] = 8'h00;
    ff_ram[4688] = 8'h00;
    ff_ram[4689] = 8'h00;
    ff_ram[4690] = 8'h00;
    ff_ram[4691] = 8'h00;
    ff_ram[4692] = 8'h00;
    ff_ram[4693] = 8'h00;
    ff_ram[4694] = 8'h00;
    ff_ram[4695] = 8'h00;
    ff_ram[4696] = 8'h00;
    ff_ram[4697] = 8'h00;
    ff_ram[4698] = 8'h00;
    ff_ram[4699] = 8'h00;
    ff_ram[4700] = 8'h00;
    ff_ram[4701] = 8'h00;
    ff_ram[4702] = 8'h00;
    ff_ram[4703] = 8'h00;
    ff_ram[4704] = 8'h00;
    ff_ram[4705] = 8'h00;
    ff_ram[4706] = 8'h00;
    ff_ram[4707] = 8'h00;
    ff_ram[4708] = 8'h00;
    ff_ram[4709] = 8'h00;
    ff_ram[4710] = 8'h00;
    ff_ram[4711] = 8'h00;
    ff_ram[4712] = 8'h00;
    ff_ram[4713] = 8'h00;
    ff_ram[4714] = 8'h00;
    ff_ram[4715] = 8'h00;
    ff_ram[4716] = 8'h00;
    ff_ram[4717] = 8'h00;
    ff_ram[4718] = 8'h00;
    ff_ram[4719] = 8'h00;
    ff_ram[4720] = 8'h00;
    ff_ram[4721] = 8'h00;
    ff_ram[4722] = 8'h00;
    ff_ram[4723] = 8'h00;
    ff_ram[4724] = 8'h00;
    ff_ram[4725] = 8'h00;
    ff_ram[4726] = 8'h00;
    ff_ram[4727] = 8'h00;
    ff_ram[4728] = 8'h00;
    ff_ram[4729] = 8'h00;
    ff_ram[4730] = 8'h00;
    ff_ram[4731] = 8'h00;
    ff_ram[4732] = 8'h00;
    ff_ram[4733] = 8'h00;
    ff_ram[4734] = 8'h00;
    ff_ram[4735] = 8'h00;
    ff_ram[4736] = 8'h00;
    ff_ram[4737] = 8'h00;
    ff_ram[4738] = 8'h00;
    ff_ram[4739] = 8'h00;
    ff_ram[4740] = 8'h00;
    ff_ram[4741] = 8'h00;
    ff_ram[4742] = 8'h00;
    ff_ram[4743] = 8'h00;
    ff_ram[4744] = 8'h00;
    ff_ram[4745] = 8'h00;
    ff_ram[4746] = 8'h00;
    ff_ram[4747] = 8'h00;
    ff_ram[4748] = 8'h00;
    ff_ram[4749] = 8'h00;
    ff_ram[4750] = 8'h00;
    ff_ram[4751] = 8'h00;
    ff_ram[4752] = 8'h00;
    ff_ram[4753] = 8'h00;
    ff_ram[4754] = 8'h00;
    ff_ram[4755] = 8'h00;
    ff_ram[4756] = 8'h00;
    ff_ram[4757] = 8'h00;
    ff_ram[4758] = 8'h00;
    ff_ram[4759] = 8'h00;
    ff_ram[4760] = 8'h00;
    ff_ram[4761] = 8'h00;
    ff_ram[4762] = 8'h00;
    ff_ram[4763] = 8'h00;
    ff_ram[4764] = 8'h00;
    ff_ram[4765] = 8'h00;
    ff_ram[4766] = 8'h00;
    ff_ram[4767] = 8'h00;
    ff_ram[4768] = 8'h00;
    ff_ram[4769] = 8'h00;
    ff_ram[4770] = 8'h00;
    ff_ram[4771] = 8'h00;
    ff_ram[4772] = 8'h00;
    ff_ram[4773] = 8'h00;
    ff_ram[4774] = 8'h00;
    ff_ram[4775] = 8'h00;
    ff_ram[4776] = 8'h00;
    ff_ram[4777] = 8'h00;
    ff_ram[4778] = 8'h00;
    ff_ram[4779] = 8'h00;
    ff_ram[4780] = 8'h00;
    ff_ram[4781] = 8'h00;
    ff_ram[4782] = 8'h00;
    ff_ram[4783] = 8'h00;
    ff_ram[4784] = 8'h00;
    ff_ram[4785] = 8'h00;
    ff_ram[4786] = 8'h00;
    ff_ram[4787] = 8'h00;
    ff_ram[4788] = 8'h00;
    ff_ram[4789] = 8'h00;
    ff_ram[4790] = 8'h00;
    ff_ram[4791] = 8'h00;
    ff_ram[4792] = 8'h00;
    ff_ram[4793] = 8'h00;
    ff_ram[4794] = 8'h00;
    ff_ram[4795] = 8'h00;
    ff_ram[4796] = 8'h00;
    ff_ram[4797] = 8'h00;
    ff_ram[4798] = 8'h00;
    ff_ram[4799] = 8'h00;
    ff_ram[4800] = 8'h00;
    ff_ram[4801] = 8'h00;
    ff_ram[4802] = 8'h00;
    ff_ram[4803] = 8'h00;
    ff_ram[4804] = 8'h00;
    ff_ram[4805] = 8'h00;
    ff_ram[4806] = 8'h00;
    ff_ram[4807] = 8'h00;
    ff_ram[4808] = 8'h00;
    ff_ram[4809] = 8'h00;
    ff_ram[4810] = 8'h00;
    ff_ram[4811] = 8'h00;
    ff_ram[4812] = 8'h00;
    ff_ram[4813] = 8'h00;
    ff_ram[4814] = 8'h00;
    ff_ram[4815] = 8'h00;
    ff_ram[4816] = 8'h00;
    ff_ram[4817] = 8'h00;
    ff_ram[4818] = 8'h00;
    ff_ram[4819] = 8'h00;
    ff_ram[4820] = 8'h00;
    ff_ram[4821] = 8'h00;
    ff_ram[4822] = 8'h00;
    ff_ram[4823] = 8'h00;
    ff_ram[4824] = 8'h00;
    ff_ram[4825] = 8'h00;
    ff_ram[4826] = 8'h00;
    ff_ram[4827] = 8'h00;
    ff_ram[4828] = 8'h00;
    ff_ram[4829] = 8'h00;
    ff_ram[4830] = 8'h00;
    ff_ram[4831] = 8'h00;
    ff_ram[4832] = 8'h00;
    ff_ram[4833] = 8'h00;
    ff_ram[4834] = 8'h00;
    ff_ram[4835] = 8'h00;
    ff_ram[4836] = 8'h00;
    ff_ram[4837] = 8'h00;
    ff_ram[4838] = 8'h00;
    ff_ram[4839] = 8'h00;
    ff_ram[4840] = 8'h00;
    ff_ram[4841] = 8'h00;
    ff_ram[4842] = 8'h00;
    ff_ram[4843] = 8'h00;
    ff_ram[4844] = 8'h00;
    ff_ram[4845] = 8'h00;
    ff_ram[4846] = 8'h00;
    ff_ram[4847] = 8'h00;
    ff_ram[4848] = 8'h00;
    ff_ram[4849] = 8'h00;
    ff_ram[4850] = 8'h00;
    ff_ram[4851] = 8'h00;
    ff_ram[4852] = 8'h00;
    ff_ram[4853] = 8'h00;
    ff_ram[4854] = 8'h00;
    ff_ram[4855] = 8'h00;
    ff_ram[4856] = 8'h00;
    ff_ram[4857] = 8'h00;
    ff_ram[4858] = 8'h00;
    ff_ram[4859] = 8'h00;
    ff_ram[4860] = 8'h00;
    ff_ram[4861] = 8'h00;
    ff_ram[4862] = 8'h00;
    ff_ram[4863] = 8'h00;
    ff_ram[4864] = 8'h00;
    ff_ram[4865] = 8'h00;
    ff_ram[4866] = 8'h00;
    ff_ram[4867] = 8'h00;
    ff_ram[4868] = 8'h00;
    ff_ram[4869] = 8'h00;
    ff_ram[4870] = 8'h00;
    ff_ram[4871] = 8'h00;
    ff_ram[4872] = 8'h00;
    ff_ram[4873] = 8'h00;
    ff_ram[4874] = 8'h00;
    ff_ram[4875] = 8'h00;
    ff_ram[4876] = 8'h00;
    ff_ram[4877] = 8'h00;
    ff_ram[4878] = 8'h00;
    ff_ram[4879] = 8'h00;
    ff_ram[4880] = 8'h00;
    ff_ram[4881] = 8'h00;
    ff_ram[4882] = 8'h00;
    ff_ram[4883] = 8'h00;
    ff_ram[4884] = 8'h00;
    ff_ram[4885] = 8'h00;
    ff_ram[4886] = 8'h00;
    ff_ram[4887] = 8'h00;
    ff_ram[4888] = 8'h00;
    ff_ram[4889] = 8'h00;
    ff_ram[4890] = 8'h00;
    ff_ram[4891] = 8'h00;
    ff_ram[4892] = 8'h00;
    ff_ram[4893] = 8'h00;
    ff_ram[4894] = 8'h00;
    ff_ram[4895] = 8'h00;
    ff_ram[4896] = 8'h00;
    ff_ram[4897] = 8'h00;
    ff_ram[4898] = 8'h00;
    ff_ram[4899] = 8'h00;
    ff_ram[4900] = 8'h00;
    ff_ram[4901] = 8'h00;
    ff_ram[4902] = 8'h00;
    ff_ram[4903] = 8'h00;
    ff_ram[4904] = 8'h00;
    ff_ram[4905] = 8'h00;
    ff_ram[4906] = 8'h00;
    ff_ram[4907] = 8'h00;
    ff_ram[4908] = 8'h00;
    ff_ram[4909] = 8'h00;
    ff_ram[4910] = 8'h00;
    ff_ram[4911] = 8'h00;
    ff_ram[4912] = 8'h00;
    ff_ram[4913] = 8'h00;
    ff_ram[4914] = 8'h00;
    ff_ram[4915] = 8'h00;
    ff_ram[4916] = 8'h00;
    ff_ram[4917] = 8'h00;
    ff_ram[4918] = 8'h00;
    ff_ram[4919] = 8'h00;
    ff_ram[4920] = 8'h00;
    ff_ram[4921] = 8'h00;
    ff_ram[4922] = 8'h00;
    ff_ram[4923] = 8'h00;
    ff_ram[4924] = 8'h00;
    ff_ram[4925] = 8'h00;
    ff_ram[4926] = 8'h00;
    ff_ram[4927] = 8'h00;
    ff_ram[4928] = 8'h00;
    ff_ram[4929] = 8'h00;
    ff_ram[4930] = 8'h00;
    ff_ram[4931] = 8'h00;
    ff_ram[4932] = 8'h00;
    ff_ram[4933] = 8'h00;
    ff_ram[4934] = 8'h00;
    ff_ram[4935] = 8'h00;
    ff_ram[4936] = 8'h00;
    ff_ram[4937] = 8'h00;
    ff_ram[4938] = 8'h00;
    ff_ram[4939] = 8'h00;
    ff_ram[4940] = 8'h00;
    ff_ram[4941] = 8'h00;
    ff_ram[4942] = 8'h00;
    ff_ram[4943] = 8'h00;
    ff_ram[4944] = 8'h00;
    ff_ram[4945] = 8'h00;
    ff_ram[4946] = 8'h00;
    ff_ram[4947] = 8'h00;
    ff_ram[4948] = 8'h00;
    ff_ram[4949] = 8'h00;
    ff_ram[4950] = 8'h00;
    ff_ram[4951] = 8'h00;
    ff_ram[4952] = 8'h00;
    ff_ram[4953] = 8'h00;
    ff_ram[4954] = 8'h00;
    ff_ram[4955] = 8'h00;
    ff_ram[4956] = 8'h00;
    ff_ram[4957] = 8'h00;
    ff_ram[4958] = 8'h00;
    ff_ram[4959] = 8'h00;
    ff_ram[4960] = 8'h00;
    ff_ram[4961] = 8'h00;
    ff_ram[4962] = 8'h00;
    ff_ram[4963] = 8'h00;
    ff_ram[4964] = 8'h00;
    ff_ram[4965] = 8'h00;
    ff_ram[4966] = 8'h00;
    ff_ram[4967] = 8'h00;
    ff_ram[4968] = 8'h00;
    ff_ram[4969] = 8'h00;
    ff_ram[4970] = 8'h00;
    ff_ram[4971] = 8'h00;
    ff_ram[4972] = 8'h00;
    ff_ram[4973] = 8'h00;
    ff_ram[4974] = 8'h00;
    ff_ram[4975] = 8'h00;
    ff_ram[4976] = 8'h00;
    ff_ram[4977] = 8'h00;
    ff_ram[4978] = 8'h00;
    ff_ram[4979] = 8'h00;
    ff_ram[4980] = 8'h00;
    ff_ram[4981] = 8'h00;
    ff_ram[4982] = 8'h00;
    ff_ram[4983] = 8'h00;
    ff_ram[4984] = 8'h00;
    ff_ram[4985] = 8'h00;
    ff_ram[4986] = 8'h00;
    ff_ram[4987] = 8'h00;
    ff_ram[4988] = 8'h00;
    ff_ram[4989] = 8'h00;
    ff_ram[4990] = 8'h00;
    ff_ram[4991] = 8'h00;
    ff_ram[4992] = 8'h00;
    ff_ram[4993] = 8'h00;
    ff_ram[4994] = 8'h00;
    ff_ram[4995] = 8'h00;
    ff_ram[4996] = 8'h00;
    ff_ram[4997] = 8'h00;
    ff_ram[4998] = 8'h00;
    ff_ram[4999] = 8'h00;
    ff_ram[5000] = 8'h00;
    ff_ram[5001] = 8'h00;
    ff_ram[5002] = 8'h00;
    ff_ram[5003] = 8'h00;
    ff_ram[5004] = 8'h00;
    ff_ram[5005] = 8'h00;
    ff_ram[5006] = 8'h00;
    ff_ram[5007] = 8'h00;
    ff_ram[5008] = 8'h00;
    ff_ram[5009] = 8'h00;
    ff_ram[5010] = 8'h00;
    ff_ram[5011] = 8'h00;
    ff_ram[5012] = 8'h00;
    ff_ram[5013] = 8'h00;
    ff_ram[5014] = 8'h00;
    ff_ram[5015] = 8'h00;
    ff_ram[5016] = 8'h00;
    ff_ram[5017] = 8'h00;
    ff_ram[5018] = 8'h00;
    ff_ram[5019] = 8'h00;
    ff_ram[5020] = 8'h00;
    ff_ram[5021] = 8'h00;
    ff_ram[5022] = 8'h00;
    ff_ram[5023] = 8'h00;
    ff_ram[5024] = 8'h00;
    ff_ram[5025] = 8'h00;
    ff_ram[5026] = 8'h00;
    ff_ram[5027] = 8'h00;
    ff_ram[5028] = 8'h00;
    ff_ram[5029] = 8'h00;
    ff_ram[5030] = 8'h00;
    ff_ram[5031] = 8'h00;
    ff_ram[5032] = 8'h00;
    ff_ram[5033] = 8'h00;
    ff_ram[5034] = 8'h00;
    ff_ram[5035] = 8'h00;
    ff_ram[5036] = 8'h00;
    ff_ram[5037] = 8'h00;
    ff_ram[5038] = 8'h00;
    ff_ram[5039] = 8'h00;
    ff_ram[5040] = 8'h00;
    ff_ram[5041] = 8'h00;
    ff_ram[5042] = 8'h00;
    ff_ram[5043] = 8'h00;
    ff_ram[5044] = 8'h00;
    ff_ram[5045] = 8'h00;
    ff_ram[5046] = 8'h00;
    ff_ram[5047] = 8'h00;
    ff_ram[5048] = 8'h00;
    ff_ram[5049] = 8'h00;
    ff_ram[5050] = 8'h00;
    ff_ram[5051] = 8'h00;
    ff_ram[5052] = 8'h00;
    ff_ram[5053] = 8'h00;
    ff_ram[5054] = 8'h00;
    ff_ram[5055] = 8'h00;
    ff_ram[5056] = 8'h00;
    ff_ram[5057] = 8'h00;
    ff_ram[5058] = 8'h00;
    ff_ram[5059] = 8'h00;
    ff_ram[5060] = 8'h00;
    ff_ram[5061] = 8'h00;
    ff_ram[5062] = 8'h00;
    ff_ram[5063] = 8'h00;
    ff_ram[5064] = 8'h00;
    ff_ram[5065] = 8'h00;
    ff_ram[5066] = 8'h00;
    ff_ram[5067] = 8'h00;
    ff_ram[5068] = 8'h00;
    ff_ram[5069] = 8'h00;
    ff_ram[5070] = 8'h00;
    ff_ram[5071] = 8'h00;
    ff_ram[5072] = 8'h00;
    ff_ram[5073] = 8'h00;
    ff_ram[5074] = 8'h00;
    ff_ram[5075] = 8'h00;
    ff_ram[5076] = 8'h00;
    ff_ram[5077] = 8'h00;
    ff_ram[5078] = 8'h00;
    ff_ram[5079] = 8'h00;
    ff_ram[5080] = 8'h00;
    ff_ram[5081] = 8'h00;
    ff_ram[5082] = 8'h00;
    ff_ram[5083] = 8'h00;
    ff_ram[5084] = 8'h00;
    ff_ram[5085] = 8'h00;
    ff_ram[5086] = 8'h00;
    ff_ram[5087] = 8'h00;
    ff_ram[5088] = 8'h00;
    ff_ram[5089] = 8'h00;
    ff_ram[5090] = 8'h00;
    ff_ram[5091] = 8'h00;
    ff_ram[5092] = 8'h00;
    ff_ram[5093] = 8'h00;
    ff_ram[5094] = 8'h00;
    ff_ram[5095] = 8'h00;
    ff_ram[5096] = 8'h00;
    ff_ram[5097] = 8'h00;
    ff_ram[5098] = 8'h00;
    ff_ram[5099] = 8'h00;
    ff_ram[5100] = 8'h00;
    ff_ram[5101] = 8'h00;
    ff_ram[5102] = 8'h00;
    ff_ram[5103] = 8'h00;
    ff_ram[5104] = 8'h00;
    ff_ram[5105] = 8'h00;
    ff_ram[5106] = 8'h00;
    ff_ram[5107] = 8'h00;
    ff_ram[5108] = 8'h00;
    ff_ram[5109] = 8'h00;
    ff_ram[5110] = 8'h00;
    ff_ram[5111] = 8'h00;
    ff_ram[5112] = 8'h00;
    ff_ram[5113] = 8'h00;
    ff_ram[5114] = 8'h00;
    ff_ram[5115] = 8'h00;
    ff_ram[5116] = 8'h00;
    ff_ram[5117] = 8'h00;
    ff_ram[5118] = 8'h00;
    ff_ram[5119] = 8'h00;
    ff_ram[5120] = 8'h00;
    ff_ram[5121] = 8'h00;
    ff_ram[5122] = 8'h00;
    ff_ram[5123] = 8'h00;
    ff_ram[5124] = 8'h00;
    ff_ram[5125] = 8'h00;
    ff_ram[5126] = 8'h00;
    ff_ram[5127] = 8'h00;
    ff_ram[5128] = 8'h00;
    ff_ram[5129] = 8'h00;
    ff_ram[5130] = 8'h00;
    ff_ram[5131] = 8'h00;
    ff_ram[5132] = 8'h00;
    ff_ram[5133] = 8'h00;
    ff_ram[5134] = 8'h00;
    ff_ram[5135] = 8'h00;
    ff_ram[5136] = 8'h00;
    ff_ram[5137] = 8'h00;
    ff_ram[5138] = 8'h00;
    ff_ram[5139] = 8'h00;
    ff_ram[5140] = 8'h00;
    ff_ram[5141] = 8'h00;
    ff_ram[5142] = 8'h00;
    ff_ram[5143] = 8'h00;
    ff_ram[5144] = 8'h00;
    ff_ram[5145] = 8'h00;
    ff_ram[5146] = 8'h00;
    ff_ram[5147] = 8'h00;
    ff_ram[5148] = 8'h00;
    ff_ram[5149] = 8'h00;
    ff_ram[5150] = 8'h00;
    ff_ram[5151] = 8'h00;
    ff_ram[5152] = 8'h00;
    ff_ram[5153] = 8'h00;
    ff_ram[5154] = 8'h00;
    ff_ram[5155] = 8'h00;
    ff_ram[5156] = 8'h00;
    ff_ram[5157] = 8'h00;
    ff_ram[5158] = 8'h00;
    ff_ram[5159] = 8'h00;
    ff_ram[5160] = 8'h00;
    ff_ram[5161] = 8'h00;
    ff_ram[5162] = 8'h00;
    ff_ram[5163] = 8'h00;
    ff_ram[5164] = 8'h00;
    ff_ram[5165] = 8'h00;
    ff_ram[5166] = 8'h00;
    ff_ram[5167] = 8'h00;
    ff_ram[5168] = 8'h00;
    ff_ram[5169] = 8'h00;
    ff_ram[5170] = 8'h00;
    ff_ram[5171] = 8'h00;
    ff_ram[5172] = 8'h00;
    ff_ram[5173] = 8'h00;
    ff_ram[5174] = 8'h00;
    ff_ram[5175] = 8'h00;
    ff_ram[5176] = 8'h00;
    ff_ram[5177] = 8'h00;
    ff_ram[5178] = 8'h00;
    ff_ram[5179] = 8'h00;
    ff_ram[5180] = 8'h00;
    ff_ram[5181] = 8'h00;
    ff_ram[5182] = 8'h00;
    ff_ram[5183] = 8'h00;
    ff_ram[5184] = 8'h00;
    ff_ram[5185] = 8'h00;
    ff_ram[5186] = 8'h00;
    ff_ram[5187] = 8'h00;
    ff_ram[5188] = 8'h00;
    ff_ram[5189] = 8'h00;
    ff_ram[5190] = 8'h00;
    ff_ram[5191] = 8'h00;
    ff_ram[5192] = 8'h00;
    ff_ram[5193] = 8'h00;
    ff_ram[5194] = 8'h00;
    ff_ram[5195] = 8'h00;
    ff_ram[5196] = 8'h00;
    ff_ram[5197] = 8'h00;
    ff_ram[5198] = 8'h00;
    ff_ram[5199] = 8'h00;
    ff_ram[5200] = 8'h00;
    ff_ram[5201] = 8'h00;
    ff_ram[5202] = 8'h00;
    ff_ram[5203] = 8'h00;
    ff_ram[5204] = 8'h00;
    ff_ram[5205] = 8'h00;
    ff_ram[5206] = 8'h00;
    ff_ram[5207] = 8'h00;
    ff_ram[5208] = 8'h00;
    ff_ram[5209] = 8'h00;
    ff_ram[5210] = 8'h00;
    ff_ram[5211] = 8'h00;
    ff_ram[5212] = 8'h00;
    ff_ram[5213] = 8'h00;
    ff_ram[5214] = 8'h00;
    ff_ram[5215] = 8'h00;
    ff_ram[5216] = 8'h00;
    ff_ram[5217] = 8'h00;
    ff_ram[5218] = 8'h00;
    ff_ram[5219] = 8'h00;
    ff_ram[5220] = 8'h00;
    ff_ram[5221] = 8'h00;
    ff_ram[5222] = 8'h00;
    ff_ram[5223] = 8'h00;
    ff_ram[5224] = 8'h00;
    ff_ram[5225] = 8'h00;
    ff_ram[5226] = 8'h00;
    ff_ram[5227] = 8'h00;
    ff_ram[5228] = 8'h00;
    ff_ram[5229] = 8'h00;
    ff_ram[5230] = 8'h00;
    ff_ram[5231] = 8'h00;
    ff_ram[5232] = 8'h00;
    ff_ram[5233] = 8'h00;
    ff_ram[5234] = 8'h00;
    ff_ram[5235] = 8'h00;
    ff_ram[5236] = 8'h00;
    ff_ram[5237] = 8'h00;
    ff_ram[5238] = 8'h00;
    ff_ram[5239] = 8'h00;
    ff_ram[5240] = 8'h00;
    ff_ram[5241] = 8'h00;
    ff_ram[5242] = 8'h00;
    ff_ram[5243] = 8'h00;
    ff_ram[5244] = 8'h00;
    ff_ram[5245] = 8'h00;
    ff_ram[5246] = 8'h00;
    ff_ram[5247] = 8'h00;
    ff_ram[5248] = 8'h00;
    ff_ram[5249] = 8'h00;
    ff_ram[5250] = 8'h00;
    ff_ram[5251] = 8'h00;
    ff_ram[5252] = 8'h00;
    ff_ram[5253] = 8'h00;
    ff_ram[5254] = 8'h00;
    ff_ram[5255] = 8'h00;
    ff_ram[5256] = 8'h00;
    ff_ram[5257] = 8'h00;
    ff_ram[5258] = 8'h00;
    ff_ram[5259] = 8'h00;
    ff_ram[5260] = 8'h00;
    ff_ram[5261] = 8'h00;
    ff_ram[5262] = 8'h00;
    ff_ram[5263] = 8'h00;
    ff_ram[5264] = 8'h00;
    ff_ram[5265] = 8'h00;
    ff_ram[5266] = 8'h00;
    ff_ram[5267] = 8'h00;
    ff_ram[5268] = 8'h00;
    ff_ram[5269] = 8'h00;
    ff_ram[5270] = 8'h00;
    ff_ram[5271] = 8'h00;
    ff_ram[5272] = 8'h00;
    ff_ram[5273] = 8'h00;
    ff_ram[5274] = 8'h00;
    ff_ram[5275] = 8'h00;
    ff_ram[5276] = 8'h00;
    ff_ram[5277] = 8'h00;
    ff_ram[5278] = 8'h00;
    ff_ram[5279] = 8'h00;
    ff_ram[5280] = 8'h00;
    ff_ram[5281] = 8'h00;
    ff_ram[5282] = 8'h00;
    ff_ram[5283] = 8'h00;
    ff_ram[5284] = 8'h00;
    ff_ram[5285] = 8'h00;
    ff_ram[5286] = 8'h00;
    ff_ram[5287] = 8'h00;
    ff_ram[5288] = 8'h00;
    ff_ram[5289] = 8'h00;
    ff_ram[5290] = 8'h00;
    ff_ram[5291] = 8'h00;
    ff_ram[5292] = 8'h00;
    ff_ram[5293] = 8'h00;
    ff_ram[5294] = 8'h00;
    ff_ram[5295] = 8'h00;
    ff_ram[5296] = 8'h00;
    ff_ram[5297] = 8'h00;
    ff_ram[5298] = 8'h00;
    ff_ram[5299] = 8'h00;
    ff_ram[5300] = 8'h00;
    ff_ram[5301] = 8'h00;
    ff_ram[5302] = 8'h00;
    ff_ram[5303] = 8'h00;
    ff_ram[5304] = 8'h00;
    ff_ram[5305] = 8'h00;
    ff_ram[5306] = 8'h00;
    ff_ram[5307] = 8'h00;
    ff_ram[5308] = 8'h00;
    ff_ram[5309] = 8'h00;
    ff_ram[5310] = 8'h00;
    ff_ram[5311] = 8'h00;
    ff_ram[5312] = 8'h00;
    ff_ram[5313] = 8'h00;
    ff_ram[5314] = 8'h00;
    ff_ram[5315] = 8'h00;
    ff_ram[5316] = 8'h00;
    ff_ram[5317] = 8'h00;
    ff_ram[5318] = 8'h00;
    ff_ram[5319] = 8'h00;
    ff_ram[5320] = 8'h00;
    ff_ram[5321] = 8'h00;
    ff_ram[5322] = 8'h00;
    ff_ram[5323] = 8'h00;
    ff_ram[5324] = 8'h00;
    ff_ram[5325] = 8'h00;
    ff_ram[5326] = 8'h00;
    ff_ram[5327] = 8'h00;
    ff_ram[5328] = 8'h00;
    ff_ram[5329] = 8'h00;
    ff_ram[5330] = 8'h00;
    ff_ram[5331] = 8'h00;
    ff_ram[5332] = 8'h00;
    ff_ram[5333] = 8'h00;
    ff_ram[5334] = 8'h00;
    ff_ram[5335] = 8'h00;
    ff_ram[5336] = 8'h00;
    ff_ram[5337] = 8'h00;
    ff_ram[5338] = 8'h00;
    ff_ram[5339] = 8'h00;
    ff_ram[5340] = 8'h00;
    ff_ram[5341] = 8'h00;
    ff_ram[5342] = 8'h00;
    ff_ram[5343] = 8'h00;
    ff_ram[5344] = 8'h00;
    ff_ram[5345] = 8'h00;
    ff_ram[5346] = 8'h00;
    ff_ram[5347] = 8'h00;
    ff_ram[5348] = 8'h00;
    ff_ram[5349] = 8'h00;
    ff_ram[5350] = 8'h00;
    ff_ram[5351] = 8'h00;
    ff_ram[5352] = 8'h00;
    ff_ram[5353] = 8'h00;
    ff_ram[5354] = 8'h00;
    ff_ram[5355] = 8'h00;
    ff_ram[5356] = 8'h00;
    ff_ram[5357] = 8'h00;
    ff_ram[5358] = 8'h00;
    ff_ram[5359] = 8'h00;
    ff_ram[5360] = 8'h00;
    ff_ram[5361] = 8'h00;
    ff_ram[5362] = 8'h00;
    ff_ram[5363] = 8'h00;
    ff_ram[5364] = 8'h00;
    ff_ram[5365] = 8'h00;
    ff_ram[5366] = 8'h00;
    ff_ram[5367] = 8'h00;
    ff_ram[5368] = 8'h00;
    ff_ram[5369] = 8'h00;
    ff_ram[5370] = 8'h00;
    ff_ram[5371] = 8'h00;
    ff_ram[5372] = 8'h00;
    ff_ram[5373] = 8'h00;
    ff_ram[5374] = 8'h00;
    ff_ram[5375] = 8'h00;
    ff_ram[5376] = 8'h00;
    ff_ram[5377] = 8'h00;
    ff_ram[5378] = 8'h00;
    ff_ram[5379] = 8'h00;
    ff_ram[5380] = 8'h00;
    ff_ram[5381] = 8'h00;
    ff_ram[5382] = 8'h00;
    ff_ram[5383] = 8'h00;
    ff_ram[5384] = 8'h00;
    ff_ram[5385] = 8'h00;
    ff_ram[5386] = 8'h00;
    ff_ram[5387] = 8'h00;
    ff_ram[5388] = 8'h00;
    ff_ram[5389] = 8'h00;
    ff_ram[5390] = 8'h00;
    ff_ram[5391] = 8'h00;
    ff_ram[5392] = 8'h00;
    ff_ram[5393] = 8'h00;
    ff_ram[5394] = 8'h00;
    ff_ram[5395] = 8'h00;
    ff_ram[5396] = 8'h00;
    ff_ram[5397] = 8'h00;
    ff_ram[5398] = 8'h00;
    ff_ram[5399] = 8'h00;
    ff_ram[5400] = 8'h00;
    ff_ram[5401] = 8'h00;
    ff_ram[5402] = 8'h00;
    ff_ram[5403] = 8'h00;
    ff_ram[5404] = 8'h00;
    ff_ram[5405] = 8'h00;
    ff_ram[5406] = 8'h00;
    ff_ram[5407] = 8'h00;
    ff_ram[5408] = 8'h00;
    ff_ram[5409] = 8'h00;
    ff_ram[5410] = 8'h00;
    ff_ram[5411] = 8'h00;
    ff_ram[5412] = 8'h00;
    ff_ram[5413] = 8'h00;
    ff_ram[5414] = 8'h00;
    ff_ram[5415] = 8'h00;
    ff_ram[5416] = 8'h00;
    ff_ram[5417] = 8'h00;
    ff_ram[5418] = 8'h00;
    ff_ram[5419] = 8'h00;
    ff_ram[5420] = 8'h00;
    ff_ram[5421] = 8'h00;
    ff_ram[5422] = 8'h00;
    ff_ram[5423] = 8'h00;
    ff_ram[5424] = 8'h00;
    ff_ram[5425] = 8'h00;
    ff_ram[5426] = 8'h00;
    ff_ram[5427] = 8'h00;
    ff_ram[5428] = 8'h00;
    ff_ram[5429] = 8'h00;
    ff_ram[5430] = 8'h00;
    ff_ram[5431] = 8'h00;
    ff_ram[5432] = 8'h00;
    ff_ram[5433] = 8'h00;
    ff_ram[5434] = 8'h00;
    ff_ram[5435] = 8'h00;
    ff_ram[5436] = 8'h00;
    ff_ram[5437] = 8'h00;
    ff_ram[5438] = 8'h00;
    ff_ram[5439] = 8'h00;
    ff_ram[5440] = 8'h00;
    ff_ram[5441] = 8'h00;
    ff_ram[5442] = 8'h00;
    ff_ram[5443] = 8'h00;
    ff_ram[5444] = 8'h00;
    ff_ram[5445] = 8'h00;
    ff_ram[5446] = 8'h00;
    ff_ram[5447] = 8'h00;
    ff_ram[5448] = 8'h00;
    ff_ram[5449] = 8'h00;
    ff_ram[5450] = 8'h00;
    ff_ram[5451] = 8'h00;
    ff_ram[5452] = 8'h00;
    ff_ram[5453] = 8'h00;
    ff_ram[5454] = 8'h00;
    ff_ram[5455] = 8'h00;
    ff_ram[5456] = 8'h00;
    ff_ram[5457] = 8'h00;
    ff_ram[5458] = 8'h00;
    ff_ram[5459] = 8'h00;
    ff_ram[5460] = 8'h00;
    ff_ram[5461] = 8'h00;
    ff_ram[5462] = 8'h00;
    ff_ram[5463] = 8'h00;
    ff_ram[5464] = 8'h00;
    ff_ram[5465] = 8'h00;
    ff_ram[5466] = 8'h00;
    ff_ram[5467] = 8'h00;
    ff_ram[5468] = 8'h00;
    ff_ram[5469] = 8'h00;
    ff_ram[5470] = 8'h00;
    ff_ram[5471] = 8'h00;
    ff_ram[5472] = 8'h00;
    ff_ram[5473] = 8'h00;
    ff_ram[5474] = 8'h00;
    ff_ram[5475] = 8'h00;
    ff_ram[5476] = 8'h00;
    ff_ram[5477] = 8'h00;
    ff_ram[5478] = 8'h00;
    ff_ram[5479] = 8'h00;
    ff_ram[5480] = 8'h00;
    ff_ram[5481] = 8'h00;
    ff_ram[5482] = 8'h00;
    ff_ram[5483] = 8'h00;
    ff_ram[5484] = 8'h00;
    ff_ram[5485] = 8'h00;
    ff_ram[5486] = 8'h00;
    ff_ram[5487] = 8'h00;
    ff_ram[5488] = 8'h00;
    ff_ram[5489] = 8'h00;
    ff_ram[5490] = 8'h00;
    ff_ram[5491] = 8'h00;
    ff_ram[5492] = 8'h00;
    ff_ram[5493] = 8'h00;
    ff_ram[5494] = 8'h00;
    ff_ram[5495] = 8'h00;
    ff_ram[5496] = 8'h00;
    ff_ram[5497] = 8'h00;
    ff_ram[5498] = 8'h00;
    ff_ram[5499] = 8'h00;
    ff_ram[5500] = 8'h00;
    ff_ram[5501] = 8'h00;
    ff_ram[5502] = 8'h00;
    ff_ram[5503] = 8'h00;
    ff_ram[5504] = 8'h00;
    ff_ram[5505] = 8'h00;
    ff_ram[5506] = 8'h00;
    ff_ram[5507] = 8'h00;
    ff_ram[5508] = 8'h00;
    ff_ram[5509] = 8'h00;
    ff_ram[5510] = 8'h00;
    ff_ram[5511] = 8'h00;
    ff_ram[5512] = 8'h00;
    ff_ram[5513] = 8'h00;
    ff_ram[5514] = 8'h00;
    ff_ram[5515] = 8'h00;
    ff_ram[5516] = 8'h00;
    ff_ram[5517] = 8'h00;
    ff_ram[5518] = 8'h00;
    ff_ram[5519] = 8'h00;
    ff_ram[5520] = 8'h00;
    ff_ram[5521] = 8'h00;
    ff_ram[5522] = 8'h00;
    ff_ram[5523] = 8'h00;
    ff_ram[5524] = 8'h00;
    ff_ram[5525] = 8'h00;
    ff_ram[5526] = 8'h00;
    ff_ram[5527] = 8'h00;
    ff_ram[5528] = 8'h00;
    ff_ram[5529] = 8'h00;
    ff_ram[5530] = 8'h00;
    ff_ram[5531] = 8'h00;
    ff_ram[5532] = 8'h00;
    ff_ram[5533] = 8'h00;
    ff_ram[5534] = 8'h00;
    ff_ram[5535] = 8'h00;
    ff_ram[5536] = 8'h00;
    ff_ram[5537] = 8'h00;
    ff_ram[5538] = 8'h00;
    ff_ram[5539] = 8'h00;
    ff_ram[5540] = 8'h00;
    ff_ram[5541] = 8'h00;
    ff_ram[5542] = 8'h00;
    ff_ram[5543] = 8'h00;
    ff_ram[5544] = 8'h00;
    ff_ram[5545] = 8'h00;
    ff_ram[5546] = 8'h00;
    ff_ram[5547] = 8'h00;
    ff_ram[5548] = 8'h00;
    ff_ram[5549] = 8'h00;
    ff_ram[5550] = 8'h00;
    ff_ram[5551] = 8'h00;
    ff_ram[5552] = 8'h00;
    ff_ram[5553] = 8'h00;
    ff_ram[5554] = 8'h00;
    ff_ram[5555] = 8'h00;
    ff_ram[5556] = 8'h00;
    ff_ram[5557] = 8'h00;
    ff_ram[5558] = 8'h00;
    ff_ram[5559] = 8'h00;
    ff_ram[5560] = 8'h00;
    ff_ram[5561] = 8'h00;
    ff_ram[5562] = 8'h00;
    ff_ram[5563] = 8'h00;
    ff_ram[5564] = 8'h00;
    ff_ram[5565] = 8'h00;
    ff_ram[5566] = 8'h00;
    ff_ram[5567] = 8'h00;
    ff_ram[5568] = 8'h00;
    ff_ram[5569] = 8'h00;
    ff_ram[5570] = 8'h00;
    ff_ram[5571] = 8'h00;
    ff_ram[5572] = 8'h00;
    ff_ram[5573] = 8'h00;
    ff_ram[5574] = 8'h00;
    ff_ram[5575] = 8'h00;
    ff_ram[5576] = 8'h00;
    ff_ram[5577] = 8'h00;
    ff_ram[5578] = 8'h00;
    ff_ram[5579] = 8'h00;
    ff_ram[5580] = 8'h00;
    ff_ram[5581] = 8'h00;
    ff_ram[5582] = 8'h00;
    ff_ram[5583] = 8'h00;
    ff_ram[5584] = 8'h00;
    ff_ram[5585] = 8'h00;
    ff_ram[5586] = 8'h00;
    ff_ram[5587] = 8'h00;
    ff_ram[5588] = 8'h00;
    ff_ram[5589] = 8'h00;
    ff_ram[5590] = 8'h00;
    ff_ram[5591] = 8'h00;
    ff_ram[5592] = 8'h00;
    ff_ram[5593] = 8'h00;
    ff_ram[5594] = 8'h00;
    ff_ram[5595] = 8'h00;
    ff_ram[5596] = 8'h00;
    ff_ram[5597] = 8'h00;
    ff_ram[5598] = 8'h00;
    ff_ram[5599] = 8'h00;
    ff_ram[5600] = 8'h00;
    ff_ram[5601] = 8'h00;
    ff_ram[5602] = 8'h00;
    ff_ram[5603] = 8'h00;
    ff_ram[5604] = 8'h00;
    ff_ram[5605] = 8'h00;
    ff_ram[5606] = 8'h00;
    ff_ram[5607] = 8'h00;
    ff_ram[5608] = 8'h00;
    ff_ram[5609] = 8'h00;
    ff_ram[5610] = 8'h00;
    ff_ram[5611] = 8'h00;
    ff_ram[5612] = 8'h00;
    ff_ram[5613] = 8'h00;
    ff_ram[5614] = 8'h00;
    ff_ram[5615] = 8'h00;
    ff_ram[5616] = 8'h00;
    ff_ram[5617] = 8'h00;
    ff_ram[5618] = 8'h00;
    ff_ram[5619] = 8'h00;
    ff_ram[5620] = 8'h00;
    ff_ram[5621] = 8'h00;
    ff_ram[5622] = 8'h00;
    ff_ram[5623] = 8'h00;
    ff_ram[5624] = 8'h00;
    ff_ram[5625] = 8'h00;
    ff_ram[5626] = 8'h00;
    ff_ram[5627] = 8'h00;
    ff_ram[5628] = 8'h00;
    ff_ram[5629] = 8'h00;
    ff_ram[5630] = 8'h00;
    ff_ram[5631] = 8'h00;
    ff_ram[5632] = 8'h00;
    ff_ram[5633] = 8'h00;
    ff_ram[5634] = 8'h00;
    ff_ram[5635] = 8'h00;
    ff_ram[5636] = 8'h00;
    ff_ram[5637] = 8'h00;
    ff_ram[5638] = 8'h00;
    ff_ram[5639] = 8'h00;
    ff_ram[5640] = 8'h00;
    ff_ram[5641] = 8'h00;
    ff_ram[5642] = 8'h00;
    ff_ram[5643] = 8'h00;
    ff_ram[5644] = 8'h00;
    ff_ram[5645] = 8'h00;
    ff_ram[5646] = 8'h00;
    ff_ram[5647] = 8'h00;
    ff_ram[5648] = 8'h00;
    ff_ram[5649] = 8'h00;
    ff_ram[5650] = 8'h00;
    ff_ram[5651] = 8'h00;
    ff_ram[5652] = 8'h00;
    ff_ram[5653] = 8'h00;
    ff_ram[5654] = 8'h00;
    ff_ram[5655] = 8'h00;
    ff_ram[5656] = 8'h00;
    ff_ram[5657] = 8'h00;
    ff_ram[5658] = 8'h00;
    ff_ram[5659] = 8'h00;
    ff_ram[5660] = 8'h00;
    ff_ram[5661] = 8'h00;
    ff_ram[5662] = 8'h00;
    ff_ram[5663] = 8'h00;
    ff_ram[5664] = 8'h00;
    ff_ram[5665] = 8'h00;
    ff_ram[5666] = 8'h00;
    ff_ram[5667] = 8'h00;
    ff_ram[5668] = 8'h00;
    ff_ram[5669] = 8'h00;
    ff_ram[5670] = 8'h00;
    ff_ram[5671] = 8'h00;
    ff_ram[5672] = 8'h00;
    ff_ram[5673] = 8'h00;
    ff_ram[5674] = 8'h00;
    ff_ram[5675] = 8'h00;
    ff_ram[5676] = 8'h00;
    ff_ram[5677] = 8'h00;
    ff_ram[5678] = 8'h00;
    ff_ram[5679] = 8'h00;
    ff_ram[5680] = 8'h00;
    ff_ram[5681] = 8'h00;
    ff_ram[5682] = 8'h00;
    ff_ram[5683] = 8'h00;
    ff_ram[5684] = 8'h00;
    ff_ram[5685] = 8'h00;
    ff_ram[5686] = 8'h00;
    ff_ram[5687] = 8'h00;
    ff_ram[5688] = 8'h00;
    ff_ram[5689] = 8'h00;
    ff_ram[5690] = 8'h00;
    ff_ram[5691] = 8'h00;
    ff_ram[5692] = 8'h00;
    ff_ram[5693] = 8'h00;
    ff_ram[5694] = 8'h00;
    ff_ram[5695] = 8'h00;
    ff_ram[5696] = 8'h00;
    ff_ram[5697] = 8'h00;
    ff_ram[5698] = 8'h00;
    ff_ram[5699] = 8'h00;
    ff_ram[5700] = 8'h00;
    ff_ram[5701] = 8'h00;
    ff_ram[5702] = 8'h00;
    ff_ram[5703] = 8'h00;
    ff_ram[5704] = 8'h00;
    ff_ram[5705] = 8'h00;
    ff_ram[5706] = 8'h00;
    ff_ram[5707] = 8'h00;
    ff_ram[5708] = 8'h00;
    ff_ram[5709] = 8'h00;
    ff_ram[5710] = 8'h00;
    ff_ram[5711] = 8'h00;
    ff_ram[5712] = 8'h00;
    ff_ram[5713] = 8'h00;
    ff_ram[5714] = 8'h00;
    ff_ram[5715] = 8'h00;
    ff_ram[5716] = 8'h00;
    ff_ram[5717] = 8'h00;
    ff_ram[5718] = 8'h00;
    ff_ram[5719] = 8'h00;
    ff_ram[5720] = 8'h00;
    ff_ram[5721] = 8'h00;
    ff_ram[5722] = 8'h00;
    ff_ram[5723] = 8'h00;
    ff_ram[5724] = 8'h00;
    ff_ram[5725] = 8'h00;
    ff_ram[5726] = 8'h00;
    ff_ram[5727] = 8'h00;
    ff_ram[5728] = 8'h00;
    ff_ram[5729] = 8'h00;
    ff_ram[5730] = 8'h00;
    ff_ram[5731] = 8'h00;
    ff_ram[5732] = 8'h00;
    ff_ram[5733] = 8'h00;
    ff_ram[5734] = 8'h00;
    ff_ram[5735] = 8'h00;
    ff_ram[5736] = 8'h00;
    ff_ram[5737] = 8'h00;
    ff_ram[5738] = 8'h00;
    ff_ram[5739] = 8'h00;
    ff_ram[5740] = 8'h00;
    ff_ram[5741] = 8'h00;
    ff_ram[5742] = 8'h00;
    ff_ram[5743] = 8'h00;
    ff_ram[5744] = 8'h00;
    ff_ram[5745] = 8'h00;
    ff_ram[5746] = 8'h00;
    ff_ram[5747] = 8'h00;
    ff_ram[5748] = 8'h00;
    ff_ram[5749] = 8'h00;
    ff_ram[5750] = 8'h00;
    ff_ram[5751] = 8'h00;
    ff_ram[5752] = 8'h00;
    ff_ram[5753] = 8'h00;
    ff_ram[5754] = 8'h00;
    ff_ram[5755] = 8'h00;
    ff_ram[5756] = 8'h00;
    ff_ram[5757] = 8'h00;
    ff_ram[5758] = 8'h00;
    ff_ram[5759] = 8'h00;
    ff_ram[5760] = 8'h00;
    ff_ram[5761] = 8'h00;
    ff_ram[5762] = 8'h00;
    ff_ram[5763] = 8'h00;
    ff_ram[5764] = 8'h00;
    ff_ram[5765] = 8'h00;
    ff_ram[5766] = 8'h00;
    ff_ram[5767] = 8'h00;
    ff_ram[5768] = 8'h00;
    ff_ram[5769] = 8'h00;
    ff_ram[5770] = 8'h00;
    ff_ram[5771] = 8'h00;
    ff_ram[5772] = 8'h00;
    ff_ram[5773] = 8'h00;
    ff_ram[5774] = 8'h00;
    ff_ram[5775] = 8'h00;
    ff_ram[5776] = 8'h00;
    ff_ram[5777] = 8'h00;
    ff_ram[5778] = 8'h00;
    ff_ram[5779] = 8'h00;
    ff_ram[5780] = 8'h00;
    ff_ram[5781] = 8'h00;
    ff_ram[5782] = 8'h00;
    ff_ram[5783] = 8'h00;
    ff_ram[5784] = 8'h00;
    ff_ram[5785] = 8'h00;
    ff_ram[5786] = 8'h00;
    ff_ram[5787] = 8'h00;
    ff_ram[5788] = 8'h00;
    ff_ram[5789] = 8'h00;
    ff_ram[5790] = 8'h00;
    ff_ram[5791] = 8'h00;
    ff_ram[5792] = 8'h00;
    ff_ram[5793] = 8'h00;
    ff_ram[5794] = 8'h00;
    ff_ram[5795] = 8'h00;
    ff_ram[5796] = 8'h00;
    ff_ram[5797] = 8'h00;
    ff_ram[5798] = 8'h00;
    ff_ram[5799] = 8'h00;
    ff_ram[5800] = 8'h00;
    ff_ram[5801] = 8'h00;
    ff_ram[5802] = 8'h00;
    ff_ram[5803] = 8'h00;
    ff_ram[5804] = 8'h00;
    ff_ram[5805] = 8'h00;
    ff_ram[5806] = 8'h00;
    ff_ram[5807] = 8'h00;
    ff_ram[5808] = 8'h00;
    ff_ram[5809] = 8'h00;
    ff_ram[5810] = 8'h00;
    ff_ram[5811] = 8'h00;
    ff_ram[5812] = 8'h00;
    ff_ram[5813] = 8'h00;
    ff_ram[5814] = 8'h00;
    ff_ram[5815] = 8'h00;
    ff_ram[5816] = 8'h00;
    ff_ram[5817] = 8'h00;
    ff_ram[5818] = 8'h00;
    ff_ram[5819] = 8'h00;
    ff_ram[5820] = 8'h00;
    ff_ram[5821] = 8'h00;
    ff_ram[5822] = 8'h00;
    ff_ram[5823] = 8'h00;
    ff_ram[5824] = 8'h00;
    ff_ram[5825] = 8'h00;
    ff_ram[5826] = 8'h00;
    ff_ram[5827] = 8'h00;
    ff_ram[5828] = 8'h00;
    ff_ram[5829] = 8'h00;
    ff_ram[5830] = 8'h00;
    ff_ram[5831] = 8'h00;
    ff_ram[5832] = 8'h00;
    ff_ram[5833] = 8'h00;
    ff_ram[5834] = 8'h00;
    ff_ram[5835] = 8'h00;
    ff_ram[5836] = 8'h00;
    ff_ram[5837] = 8'h00;
    ff_ram[5838] = 8'h00;
    ff_ram[5839] = 8'h00;
    ff_ram[5840] = 8'h00;
    ff_ram[5841] = 8'h00;
    ff_ram[5842] = 8'h00;
    ff_ram[5843] = 8'h00;
    ff_ram[5844] = 8'h00;
    ff_ram[5845] = 8'h00;
    ff_ram[5846] = 8'h00;
    ff_ram[5847] = 8'h00;
    ff_ram[5848] = 8'h00;
    ff_ram[5849] = 8'h00;
    ff_ram[5850] = 8'h00;
    ff_ram[5851] = 8'h00;
    ff_ram[5852] = 8'h00;
    ff_ram[5853] = 8'h00;
    ff_ram[5854] = 8'h00;
    ff_ram[5855] = 8'h00;
    ff_ram[5856] = 8'h00;
    ff_ram[5857] = 8'h00;
    ff_ram[5858] = 8'h00;
    ff_ram[5859] = 8'h00;
    ff_ram[5860] = 8'h00;
    ff_ram[5861] = 8'h00;
    ff_ram[5862] = 8'h00;
    ff_ram[5863] = 8'h00;
    ff_ram[5864] = 8'h00;
    ff_ram[5865] = 8'h00;
    ff_ram[5866] = 8'h00;
    ff_ram[5867] = 8'h00;
    ff_ram[5868] = 8'h00;
    ff_ram[5869] = 8'h00;
    ff_ram[5870] = 8'h00;
    ff_ram[5871] = 8'h00;
    ff_ram[5872] = 8'h00;
    ff_ram[5873] = 8'h00;
    ff_ram[5874] = 8'h00;
    ff_ram[5875] = 8'h00;
    ff_ram[5876] = 8'h00;
    ff_ram[5877] = 8'h00;
    ff_ram[5878] = 8'h00;
    ff_ram[5879] = 8'h00;
    ff_ram[5880] = 8'h00;
    ff_ram[5881] = 8'h00;
    ff_ram[5882] = 8'h00;
    ff_ram[5883] = 8'h00;
    ff_ram[5884] = 8'h00;
    ff_ram[5885] = 8'h00;
    ff_ram[5886] = 8'h00;
    ff_ram[5887] = 8'h00;
    ff_ram[5888] = 8'h00;
    ff_ram[5889] = 8'h00;
    ff_ram[5890] = 8'h00;
    ff_ram[5891] = 8'h00;
    ff_ram[5892] = 8'h00;
    ff_ram[5893] = 8'h00;
    ff_ram[5894] = 8'h00;
    ff_ram[5895] = 8'h00;
    ff_ram[5896] = 8'h00;
    ff_ram[5897] = 8'h00;
    ff_ram[5898] = 8'h00;
    ff_ram[5899] = 8'h00;
    ff_ram[5900] = 8'h00;
    ff_ram[5901] = 8'h00;
    ff_ram[5902] = 8'h00;
    ff_ram[5903] = 8'h00;
    ff_ram[5904] = 8'h00;
    ff_ram[5905] = 8'h00;
    ff_ram[5906] = 8'h00;
    ff_ram[5907] = 8'h00;
    ff_ram[5908] = 8'h00;
    ff_ram[5909] = 8'h00;
    ff_ram[5910] = 8'h00;
    ff_ram[5911] = 8'h00;
    ff_ram[5912] = 8'h00;
    ff_ram[5913] = 8'h00;
    ff_ram[5914] = 8'h00;
    ff_ram[5915] = 8'h00;
    ff_ram[5916] = 8'h00;
    ff_ram[5917] = 8'h00;
    ff_ram[5918] = 8'h00;
    ff_ram[5919] = 8'h00;
    ff_ram[5920] = 8'h00;
    ff_ram[5921] = 8'h00;
    ff_ram[5922] = 8'h00;
    ff_ram[5923] = 8'h00;
    ff_ram[5924] = 8'h00;
    ff_ram[5925] = 8'h00;
    ff_ram[5926] = 8'h00;
    ff_ram[5927] = 8'h00;
    ff_ram[5928] = 8'h00;
    ff_ram[5929] = 8'h00;
    ff_ram[5930] = 8'h00;
    ff_ram[5931] = 8'h00;
    ff_ram[5932] = 8'h00;
    ff_ram[5933] = 8'h00;
    ff_ram[5934] = 8'h00;
    ff_ram[5935] = 8'h00;
    ff_ram[5936] = 8'h00;
    ff_ram[5937] = 8'h00;
    ff_ram[5938] = 8'h00;
    ff_ram[5939] = 8'h00;
    ff_ram[5940] = 8'h00;
    ff_ram[5941] = 8'h00;
    ff_ram[5942] = 8'h00;
    ff_ram[5943] = 8'h00;
    ff_ram[5944] = 8'h00;
    ff_ram[5945] = 8'h00;
    ff_ram[5946] = 8'h00;
    ff_ram[5947] = 8'h00;
    ff_ram[5948] = 8'h00;
    ff_ram[5949] = 8'h00;
    ff_ram[5950] = 8'h00;
    ff_ram[5951] = 8'h00;
    ff_ram[5952] = 8'h00;
    ff_ram[5953] = 8'h00;
    ff_ram[5954] = 8'h00;
    ff_ram[5955] = 8'h00;
    ff_ram[5956] = 8'h00;
    ff_ram[5957] = 8'h00;
    ff_ram[5958] = 8'h00;
    ff_ram[5959] = 8'h00;
    ff_ram[5960] = 8'h00;
    ff_ram[5961] = 8'h00;
    ff_ram[5962] = 8'h00;
    ff_ram[5963] = 8'h00;
    ff_ram[5964] = 8'h00;
    ff_ram[5965] = 8'h00;
    ff_ram[5966] = 8'h00;
    ff_ram[5967] = 8'h00;
    ff_ram[5968] = 8'h00;
    ff_ram[5969] = 8'h00;
    ff_ram[5970] = 8'h00;
    ff_ram[5971] = 8'h00;
    ff_ram[5972] = 8'h00;
    ff_ram[5973] = 8'h00;
    ff_ram[5974] = 8'h00;
    ff_ram[5975] = 8'h00;
    ff_ram[5976] = 8'h00;
    ff_ram[5977] = 8'h00;
    ff_ram[5978] = 8'h00;
    ff_ram[5979] = 8'h00;
    ff_ram[5980] = 8'h00;
    ff_ram[5981] = 8'h00;
    ff_ram[5982] = 8'h00;
    ff_ram[5983] = 8'h00;
    ff_ram[5984] = 8'h00;
    ff_ram[5985] = 8'h00;
    ff_ram[5986] = 8'h00;
    ff_ram[5987] = 8'h00;
    ff_ram[5988] = 8'h00;
    ff_ram[5989] = 8'h00;
    ff_ram[5990] = 8'h00;
    ff_ram[5991] = 8'h00;
    ff_ram[5992] = 8'h00;
    ff_ram[5993] = 8'h00;
    ff_ram[5994] = 8'h00;
    ff_ram[5995] = 8'h00;
    ff_ram[5996] = 8'h00;
    ff_ram[5997] = 8'h00;
    ff_ram[5998] = 8'h00;
    ff_ram[5999] = 8'h00;
    ff_ram[6000] = 8'h00;
    ff_ram[6001] = 8'h00;
    ff_ram[6002] = 8'h00;
    ff_ram[6003] = 8'h00;
    ff_ram[6004] = 8'h00;
    ff_ram[6005] = 8'h00;
    ff_ram[6006] = 8'h00;
    ff_ram[6007] = 8'h00;
    ff_ram[6008] = 8'h00;
    ff_ram[6009] = 8'h00;
    ff_ram[6010] = 8'h00;
    ff_ram[6011] = 8'h00;
    ff_ram[6012] = 8'h00;
    ff_ram[6013] = 8'h00;
    ff_ram[6014] = 8'h00;
    ff_ram[6015] = 8'h00;
    ff_ram[6016] = 8'h00;
    ff_ram[6017] = 8'h00;
    ff_ram[6018] = 8'h00;
    ff_ram[6019] = 8'h00;
    ff_ram[6020] = 8'h00;
    ff_ram[6021] = 8'h00;
    ff_ram[6022] = 8'h00;
    ff_ram[6023] = 8'h00;
    ff_ram[6024] = 8'h00;
    ff_ram[6025] = 8'h00;
    ff_ram[6026] = 8'h00;
    ff_ram[6027] = 8'h00;
    ff_ram[6028] = 8'h00;
    ff_ram[6029] = 8'h00;
    ff_ram[6030] = 8'h00;
    ff_ram[6031] = 8'h00;
    ff_ram[6032] = 8'h00;
    ff_ram[6033] = 8'h00;
    ff_ram[6034] = 8'h00;
    ff_ram[6035] = 8'h00;
    ff_ram[6036] = 8'h00;
    ff_ram[6037] = 8'h00;
    ff_ram[6038] = 8'h00;
    ff_ram[6039] = 8'h00;
    ff_ram[6040] = 8'h00;
    ff_ram[6041] = 8'h00;
    ff_ram[6042] = 8'h00;
    ff_ram[6043] = 8'h00;
    ff_ram[6044] = 8'h00;
    ff_ram[6045] = 8'h00;
    ff_ram[6046] = 8'h00;
    ff_ram[6047] = 8'h00;
    ff_ram[6048] = 8'h00;
    ff_ram[6049] = 8'h00;
    ff_ram[6050] = 8'h00;
    ff_ram[6051] = 8'h00;
    ff_ram[6052] = 8'h00;
    ff_ram[6053] = 8'h00;
    ff_ram[6054] = 8'h00;
    ff_ram[6055] = 8'h00;
    ff_ram[6056] = 8'h00;
    ff_ram[6057] = 8'h00;
    ff_ram[6058] = 8'h00;
    ff_ram[6059] = 8'h00;
    ff_ram[6060] = 8'h00;
    ff_ram[6061] = 8'h00;
    ff_ram[6062] = 8'h00;
    ff_ram[6063] = 8'h00;
    ff_ram[6064] = 8'h00;
    ff_ram[6065] = 8'h00;
    ff_ram[6066] = 8'h00;
    ff_ram[6067] = 8'h00;
    ff_ram[6068] = 8'h00;
    ff_ram[6069] = 8'h00;
    ff_ram[6070] = 8'h00;
    ff_ram[6071] = 8'h00;
    ff_ram[6072] = 8'h00;
    ff_ram[6073] = 8'h00;
    ff_ram[6074] = 8'h00;
    ff_ram[6075] = 8'h00;
    ff_ram[6076] = 8'h00;
    ff_ram[6077] = 8'h00;
    ff_ram[6078] = 8'h00;
    ff_ram[6079] = 8'h00;
    ff_ram[6080] = 8'h00;
    ff_ram[6081] = 8'h00;
    ff_ram[6082] = 8'h00;
    ff_ram[6083] = 8'h00;
    ff_ram[6084] = 8'h00;
    ff_ram[6085] = 8'h00;
    ff_ram[6086] = 8'h00;
    ff_ram[6087] = 8'h00;
    ff_ram[6088] = 8'h00;
    ff_ram[6089] = 8'h00;
    ff_ram[6090] = 8'h00;
    ff_ram[6091] = 8'h00;
    ff_ram[6092] = 8'h00;
    ff_ram[6093] = 8'h00;
    ff_ram[6094] = 8'h00;
    ff_ram[6095] = 8'h00;
    ff_ram[6096] = 8'h00;
    ff_ram[6097] = 8'h00;
    ff_ram[6098] = 8'h00;
    ff_ram[6099] = 8'h00;
    ff_ram[6100] = 8'h00;
    ff_ram[6101] = 8'h00;
    ff_ram[6102] = 8'h00;
    ff_ram[6103] = 8'h00;
    ff_ram[6104] = 8'h00;
    ff_ram[6105] = 8'h00;
    ff_ram[6106] = 8'h00;
    ff_ram[6107] = 8'h00;
    ff_ram[6108] = 8'h00;
    ff_ram[6109] = 8'h00;
    ff_ram[6110] = 8'h00;
    ff_ram[6111] = 8'h00;
    ff_ram[6112] = 8'h00;
    ff_ram[6113] = 8'h00;
    ff_ram[6114] = 8'h00;
    ff_ram[6115] = 8'h00;
    ff_ram[6116] = 8'h00;
    ff_ram[6117] = 8'h00;
    ff_ram[6118] = 8'h00;
    ff_ram[6119] = 8'h00;
    ff_ram[6120] = 8'h00;
    ff_ram[6121] = 8'h00;
    ff_ram[6122] = 8'h00;
    ff_ram[6123] = 8'h00;
    ff_ram[6124] = 8'h00;
    ff_ram[6125] = 8'h00;
    ff_ram[6126] = 8'h00;
    ff_ram[6127] = 8'h00;
    ff_ram[6128] = 8'h00;
    ff_ram[6129] = 8'h00;
    ff_ram[6130] = 8'h00;
    ff_ram[6131] = 8'h00;
    ff_ram[6132] = 8'h00;
    ff_ram[6133] = 8'h00;
    ff_ram[6134] = 8'h00;
    ff_ram[6135] = 8'h00;
    ff_ram[6136] = 8'h00;
    ff_ram[6137] = 8'h00;
    ff_ram[6138] = 8'h00;
    ff_ram[6139] = 8'h00;
    ff_ram[6140] = 8'h00;
    ff_ram[6141] = 8'h00;
    ff_ram[6142] = 8'h00;
    ff_ram[6143] = 8'h00;
    ff_ram[6144] = 8'h20;
    ff_ram[6145] = 8'h20;
    ff_ram[6146] = 8'h4D;
    ff_ram[6147] = 8'h53;
    ff_ram[6148] = 8'h58;
    ff_ram[6149] = 8'h20;
    ff_ram[6150] = 8'h42;
    ff_ram[6151] = 8'h41;
    ff_ram[6152] = 8'h53;
    ff_ram[6153] = 8'h49;
    ff_ram[6154] = 8'h43;
    ff_ram[6155] = 8'h20;
    ff_ram[6156] = 8'h76;
    ff_ram[6157] = 8'h65;
    ff_ram[6158] = 8'h72;
    ff_ram[6159] = 8'h73;
    ff_ram[6160] = 8'h69;
    ff_ram[6161] = 8'h6F;
    ff_ram[6162] = 8'h6E;
    ff_ram[6163] = 8'h20;
    ff_ram[6164] = 8'h34;
    ff_ram[6165] = 8'h2E;
    ff_ram[6166] = 8'h31;
    ff_ram[6167] = 8'h20;
    ff_ram[6168] = 8'h20;
    ff_ram[6169] = 8'h20;
    ff_ram[6170] = 8'h20;
    ff_ram[6171] = 8'h20;
    ff_ram[6172] = 8'h20;
    ff_ram[6173] = 8'h20;
    ff_ram[6174] = 8'h20;
    ff_ram[6175] = 8'h20;
    ff_ram[6176] = 8'h20;
    ff_ram[6177] = 8'h20;
    ff_ram[6178] = 8'h43;
    ff_ram[6179] = 8'h6F;
    ff_ram[6180] = 8'h70;
    ff_ram[6181] = 8'h79;
    ff_ram[6182] = 8'h72;
    ff_ram[6183] = 8'h69;
    ff_ram[6184] = 8'h67;
    ff_ram[6185] = 8'h68;
    ff_ram[6186] = 8'h74;
    ff_ram[6187] = 8'h20;
    ff_ram[6188] = 8'h31;
    ff_ram[6189] = 8'h39;
    ff_ram[6190] = 8'h39;
    ff_ram[6191] = 8'h30;
    ff_ram[6192] = 8'h20;
    ff_ram[6193] = 8'h62;
    ff_ram[6194] = 8'h79;
    ff_ram[6195] = 8'h20;
    ff_ram[6196] = 8'h4D;
    ff_ram[6197] = 8'h69;
    ff_ram[6198] = 8'h63;
    ff_ram[6199] = 8'h72;
    ff_ram[6200] = 8'h6F;
    ff_ram[6201] = 8'h73;
    ff_ram[6202] = 8'h6F;
    ff_ram[6203] = 8'h66;
    ff_ram[6204] = 8'h74;
    ff_ram[6205] = 8'h20;
    ff_ram[6206] = 8'h20;
    ff_ram[6207] = 8'h20;
    ff_ram[6208] = 8'h20;
    ff_ram[6209] = 8'h20;
    ff_ram[6210] = 8'h32;
    ff_ram[6211] = 8'h35;
    ff_ram[6212] = 8'h32;
    ff_ram[6213] = 8'h37;
    ff_ram[6214] = 8'h31;
    ff_ram[6215] = 8'h20;
    ff_ram[6216] = 8'h42;
    ff_ram[6217] = 8'h79;
    ff_ram[6218] = 8'h74;
    ff_ram[6219] = 8'h65;
    ff_ram[6220] = 8'h73;
    ff_ram[6221] = 8'h20;
    ff_ram[6222] = 8'h66;
    ff_ram[6223] = 8'h72;
    ff_ram[6224] = 8'h65;
    ff_ram[6225] = 8'h65;
    ff_ram[6226] = 8'h20;
    ff_ram[6227] = 8'h20;
    ff_ram[6228] = 8'h20;
    ff_ram[6229] = 8'h20;
    ff_ram[6230] = 8'h20;
    ff_ram[6231] = 8'h20;
    ff_ram[6232] = 8'h20;
    ff_ram[6233] = 8'h20;
    ff_ram[6234] = 8'h20;
    ff_ram[6235] = 8'h20;
    ff_ram[6236] = 8'h20;
    ff_ram[6237] = 8'h20;
    ff_ram[6238] = 8'h20;
    ff_ram[6239] = 8'h20;
    ff_ram[6240] = 8'h20;
    ff_ram[6241] = 8'h20;
    ff_ram[6242] = 8'h44;
    ff_ram[6243] = 8'h69;
    ff_ram[6244] = 8'h73;
    ff_ram[6245] = 8'h6B;
    ff_ram[6246] = 8'h20;
    ff_ram[6247] = 8'h42;
    ff_ram[6248] = 8'h41;
    ff_ram[6249] = 8'h53;
    ff_ram[6250] = 8'h49;
    ff_ram[6251] = 8'h43;
    ff_ram[6252] = 8'h20;
    ff_ram[6253] = 8'h76;
    ff_ram[6254] = 8'h65;
    ff_ram[6255] = 8'h72;
    ff_ram[6256] = 8'h73;
    ff_ram[6257] = 8'h69;
    ff_ram[6258] = 8'h6F;
    ff_ram[6259] = 8'h6E;
    ff_ram[6260] = 8'h20;
    ff_ram[6261] = 8'h32;
    ff_ram[6262] = 8'h2E;
    ff_ram[6263] = 8'h30;
    ff_ram[6264] = 8'h31;
    ff_ram[6265] = 8'h20;
    ff_ram[6266] = 8'h20;
    ff_ram[6267] = 8'h20;
    ff_ram[6268] = 8'h20;
    ff_ram[6269] = 8'h20;
    ff_ram[6270] = 8'h20;
    ff_ram[6271] = 8'h20;
    ff_ram[6272] = 8'h20;
    ff_ram[6273] = 8'h20;
    ff_ram[6274] = 8'h4F;
    ff_ram[6275] = 8'h6B;
    ff_ram[6276] = 8'h20;
    ff_ram[6277] = 8'h20;
    ff_ram[6278] = 8'h20;
    ff_ram[6279] = 8'h20;
    ff_ram[6280] = 8'h20;
    ff_ram[6281] = 8'h20;
    ff_ram[6282] = 8'h20;
    ff_ram[6283] = 8'h20;
    ff_ram[6284] = 8'h20;
    ff_ram[6285] = 8'h20;
    ff_ram[6286] = 8'h20;
    ff_ram[6287] = 8'h20;
    ff_ram[6288] = 8'h20;
    ff_ram[6289] = 8'h20;
    ff_ram[6290] = 8'h20;
    ff_ram[6291] = 8'h20;
    ff_ram[6292] = 8'h20;
    ff_ram[6293] = 8'h20;
    ff_ram[6294] = 8'h20;
    ff_ram[6295] = 8'h20;
    ff_ram[6296] = 8'h20;
    ff_ram[6297] = 8'h20;
    ff_ram[6298] = 8'h20;
    ff_ram[6299] = 8'h20;
    ff_ram[6300] = 8'h20;
    ff_ram[6301] = 8'h20;
    ff_ram[6302] = 8'h20;
    ff_ram[6303] = 8'h20;
    ff_ram[6304] = 8'h20;
    ff_ram[6305] = 8'h20;
    ff_ram[6306] = 8'h62;
    ff_ram[6307] = 8'h73;
    ff_ram[6308] = 8'h61;
    ff_ram[6309] = 8'h76;
    ff_ram[6310] = 8'h65;
    ff_ram[6311] = 8'h20;
    ff_ram[6312] = 8'h22;
    ff_ram[6313] = 8'h76;
    ff_ram[6314] = 8'h72;
    ff_ram[6315] = 8'h61;
    ff_ram[6316] = 8'h6D;
    ff_ram[6317] = 8'h2E;
    ff_ram[6318] = 8'h62;
    ff_ram[6319] = 8'h69;
    ff_ram[6320] = 8'h6E;
    ff_ram[6321] = 8'h22;
    ff_ram[6322] = 8'h2C;
    ff_ram[6323] = 8'h30;
    ff_ram[6324] = 8'h2C;
    ff_ram[6325] = 8'h26;
    ff_ram[6326] = 8'h48;
    ff_ram[6327] = 8'h33;
    ff_ram[6328] = 8'h46;
    ff_ram[6329] = 8'h46;
    ff_ram[6330] = 8'h46;
    ff_ram[6331] = 8'h2C;
    ff_ram[6332] = 8'h53;
    ff_ram[6333] = 8'h20;
    ff_ram[6334] = 8'h20;
    ff_ram[6335] = 8'h20;
    ff_ram[6336] = 8'h20;
    ff_ram[6337] = 8'h20;
    ff_ram[6338] = 8'h20;
    ff_ram[6339] = 8'h20;
    ff_ram[6340] = 8'h20;
    ff_ram[6341] = 8'h20;
    ff_ram[6342] = 8'h20;
    ff_ram[6343] = 8'h20;
    ff_ram[6344] = 8'h20;
    ff_ram[6345] = 8'h20;
    ff_ram[6346] = 8'h20;
    ff_ram[6347] = 8'h20;
    ff_ram[6348] = 8'h20;
    ff_ram[6349] = 8'h20;
    ff_ram[6350] = 8'h20;
    ff_ram[6351] = 8'h20;
    ff_ram[6352] = 8'h20;
    ff_ram[6353] = 8'h20;
    ff_ram[6354] = 8'h20;
    ff_ram[6355] = 8'h20;
    ff_ram[6356] = 8'h20;
    ff_ram[6357] = 8'h20;
    ff_ram[6358] = 8'h20;
    ff_ram[6359] = 8'h20;
    ff_ram[6360] = 8'h20;
    ff_ram[6361] = 8'h20;
    ff_ram[6362] = 8'h20;
    ff_ram[6363] = 8'h20;
    ff_ram[6364] = 8'h20;
    ff_ram[6365] = 8'h20;
    ff_ram[6366] = 8'h20;
    ff_ram[6367] = 8'h20;
    ff_ram[6368] = 8'h20;
    ff_ram[6369] = 8'h20;
    ff_ram[6370] = 8'h20;
    ff_ram[6371] = 8'h20;
    ff_ram[6372] = 8'h20;
    ff_ram[6373] = 8'h20;
    ff_ram[6374] = 8'h20;
    ff_ram[6375] = 8'h20;
    ff_ram[6376] = 8'h20;
    ff_ram[6377] = 8'h20;
    ff_ram[6378] = 8'h20;
    ff_ram[6379] = 8'h20;
    ff_ram[6380] = 8'h20;
    ff_ram[6381] = 8'h20;
    ff_ram[6382] = 8'h20;
    ff_ram[6383] = 8'h20;
    ff_ram[6384] = 8'h20;
    ff_ram[6385] = 8'h20;
    ff_ram[6386] = 8'h20;
    ff_ram[6387] = 8'h20;
    ff_ram[6388] = 8'h20;
    ff_ram[6389] = 8'h20;
    ff_ram[6390] = 8'h20;
    ff_ram[6391] = 8'h20;
    ff_ram[6392] = 8'h20;
    ff_ram[6393] = 8'h20;
    ff_ram[6394] = 8'h20;
    ff_ram[6395] = 8'h20;
    ff_ram[6396] = 8'h20;
    ff_ram[6397] = 8'h20;
    ff_ram[6398] = 8'h20;
    ff_ram[6399] = 8'h20;
    ff_ram[6400] = 8'h20;
    ff_ram[6401] = 8'h20;
    ff_ram[6402] = 8'h20;
    ff_ram[6403] = 8'h20;
    ff_ram[6404] = 8'h20;
    ff_ram[6405] = 8'h20;
    ff_ram[6406] = 8'h20;
    ff_ram[6407] = 8'h20;
    ff_ram[6408] = 8'h20;
    ff_ram[6409] = 8'h20;
    ff_ram[6410] = 8'h20;
    ff_ram[6411] = 8'h20;
    ff_ram[6412] = 8'h20;
    ff_ram[6413] = 8'h20;
    ff_ram[6414] = 8'h20;
    ff_ram[6415] = 8'h20;
    ff_ram[6416] = 8'h20;
    ff_ram[6417] = 8'h20;
    ff_ram[6418] = 8'h20;
    ff_ram[6419] = 8'h20;
    ff_ram[6420] = 8'h20;
    ff_ram[6421] = 8'h20;
    ff_ram[6422] = 8'h20;
    ff_ram[6423] = 8'h20;
    ff_ram[6424] = 8'h20;
    ff_ram[6425] = 8'h20;
    ff_ram[6426] = 8'h20;
    ff_ram[6427] = 8'h20;
    ff_ram[6428] = 8'h20;
    ff_ram[6429] = 8'h20;
    ff_ram[6430] = 8'h20;
    ff_ram[6431] = 8'h20;
    ff_ram[6432] = 8'h20;
    ff_ram[6433] = 8'h20;
    ff_ram[6434] = 8'h20;
    ff_ram[6435] = 8'h20;
    ff_ram[6436] = 8'h20;
    ff_ram[6437] = 8'h20;
    ff_ram[6438] = 8'h20;
    ff_ram[6439] = 8'h20;
    ff_ram[6440] = 8'h20;
    ff_ram[6441] = 8'h20;
    ff_ram[6442] = 8'h20;
    ff_ram[6443] = 8'h20;
    ff_ram[6444] = 8'h20;
    ff_ram[6445] = 8'h20;
    ff_ram[6446] = 8'h20;
    ff_ram[6447] = 8'h20;
    ff_ram[6448] = 8'h20;
    ff_ram[6449] = 8'h20;
    ff_ram[6450] = 8'h20;
    ff_ram[6451] = 8'h20;
    ff_ram[6452] = 8'h20;
    ff_ram[6453] = 8'h20;
    ff_ram[6454] = 8'h20;
    ff_ram[6455] = 8'h20;
    ff_ram[6456] = 8'h20;
    ff_ram[6457] = 8'h20;
    ff_ram[6458] = 8'h20;
    ff_ram[6459] = 8'h20;
    ff_ram[6460] = 8'h20;
    ff_ram[6461] = 8'h20;
    ff_ram[6462] = 8'h20;
    ff_ram[6463] = 8'h20;
    ff_ram[6464] = 8'h20;
    ff_ram[6465] = 8'h20;
    ff_ram[6466] = 8'h20;
    ff_ram[6467] = 8'h20;
    ff_ram[6468] = 8'h20;
    ff_ram[6469] = 8'h20;
    ff_ram[6470] = 8'h20;
    ff_ram[6471] = 8'h20;
    ff_ram[6472] = 8'h20;
    ff_ram[6473] = 8'h20;
    ff_ram[6474] = 8'h20;
    ff_ram[6475] = 8'h20;
    ff_ram[6476] = 8'h20;
    ff_ram[6477] = 8'h20;
    ff_ram[6478] = 8'h20;
    ff_ram[6479] = 8'h20;
    ff_ram[6480] = 8'h20;
    ff_ram[6481] = 8'h20;
    ff_ram[6482] = 8'h20;
    ff_ram[6483] = 8'h20;
    ff_ram[6484] = 8'h20;
    ff_ram[6485] = 8'h20;
    ff_ram[6486] = 8'h20;
    ff_ram[6487] = 8'h20;
    ff_ram[6488] = 8'h20;
    ff_ram[6489] = 8'h20;
    ff_ram[6490] = 8'h20;
    ff_ram[6491] = 8'h20;
    ff_ram[6492] = 8'h20;
    ff_ram[6493] = 8'h20;
    ff_ram[6494] = 8'h20;
    ff_ram[6495] = 8'h20;
    ff_ram[6496] = 8'h20;
    ff_ram[6497] = 8'h20;
    ff_ram[6498] = 8'h20;
    ff_ram[6499] = 8'h20;
    ff_ram[6500] = 8'h20;
    ff_ram[6501] = 8'h20;
    ff_ram[6502] = 8'h20;
    ff_ram[6503] = 8'h20;
    ff_ram[6504] = 8'h20;
    ff_ram[6505] = 8'h20;
    ff_ram[6506] = 8'h20;
    ff_ram[6507] = 8'h20;
    ff_ram[6508] = 8'h20;
    ff_ram[6509] = 8'h20;
    ff_ram[6510] = 8'h20;
    ff_ram[6511] = 8'h20;
    ff_ram[6512] = 8'h20;
    ff_ram[6513] = 8'h20;
    ff_ram[6514] = 8'h20;
    ff_ram[6515] = 8'h20;
    ff_ram[6516] = 8'h20;
    ff_ram[6517] = 8'h20;
    ff_ram[6518] = 8'h20;
    ff_ram[6519] = 8'h20;
    ff_ram[6520] = 8'h20;
    ff_ram[6521] = 8'h20;
    ff_ram[6522] = 8'h20;
    ff_ram[6523] = 8'h20;
    ff_ram[6524] = 8'h20;
    ff_ram[6525] = 8'h20;
    ff_ram[6526] = 8'h20;
    ff_ram[6527] = 8'h20;
    ff_ram[6528] = 8'h20;
    ff_ram[6529] = 8'h20;
    ff_ram[6530] = 8'h20;
    ff_ram[6531] = 8'h20;
    ff_ram[6532] = 8'h20;
    ff_ram[6533] = 8'h20;
    ff_ram[6534] = 8'h20;
    ff_ram[6535] = 8'h20;
    ff_ram[6536] = 8'h20;
    ff_ram[6537] = 8'h20;
    ff_ram[6538] = 8'h20;
    ff_ram[6539] = 8'h20;
    ff_ram[6540] = 8'h20;
    ff_ram[6541] = 8'h20;
    ff_ram[6542] = 8'h20;
    ff_ram[6543] = 8'h20;
    ff_ram[6544] = 8'h20;
    ff_ram[6545] = 8'h20;
    ff_ram[6546] = 8'h20;
    ff_ram[6547] = 8'h20;
    ff_ram[6548] = 8'h20;
    ff_ram[6549] = 8'h20;
    ff_ram[6550] = 8'h20;
    ff_ram[6551] = 8'h20;
    ff_ram[6552] = 8'h20;
    ff_ram[6553] = 8'h20;
    ff_ram[6554] = 8'h20;
    ff_ram[6555] = 8'h20;
    ff_ram[6556] = 8'h20;
    ff_ram[6557] = 8'h20;
    ff_ram[6558] = 8'h20;
    ff_ram[6559] = 8'h20;
    ff_ram[6560] = 8'h20;
    ff_ram[6561] = 8'h20;
    ff_ram[6562] = 8'h20;
    ff_ram[6563] = 8'h20;
    ff_ram[6564] = 8'h20;
    ff_ram[6565] = 8'h20;
    ff_ram[6566] = 8'h20;
    ff_ram[6567] = 8'h20;
    ff_ram[6568] = 8'h20;
    ff_ram[6569] = 8'h20;
    ff_ram[6570] = 8'h20;
    ff_ram[6571] = 8'h20;
    ff_ram[6572] = 8'h20;
    ff_ram[6573] = 8'h20;
    ff_ram[6574] = 8'h20;
    ff_ram[6575] = 8'h20;
    ff_ram[6576] = 8'h20;
    ff_ram[6577] = 8'h20;
    ff_ram[6578] = 8'h20;
    ff_ram[6579] = 8'h20;
    ff_ram[6580] = 8'h20;
    ff_ram[6581] = 8'h20;
    ff_ram[6582] = 8'h20;
    ff_ram[6583] = 8'h20;
    ff_ram[6584] = 8'h20;
    ff_ram[6585] = 8'h20;
    ff_ram[6586] = 8'h20;
    ff_ram[6587] = 8'h20;
    ff_ram[6588] = 8'h20;
    ff_ram[6589] = 8'h20;
    ff_ram[6590] = 8'h20;
    ff_ram[6591] = 8'h20;
    ff_ram[6592] = 8'h20;
    ff_ram[6593] = 8'h20;
    ff_ram[6594] = 8'h20;
    ff_ram[6595] = 8'h20;
    ff_ram[6596] = 8'h20;
    ff_ram[6597] = 8'h20;
    ff_ram[6598] = 8'h20;
    ff_ram[6599] = 8'h20;
    ff_ram[6600] = 8'h20;
    ff_ram[6601] = 8'h20;
    ff_ram[6602] = 8'h20;
    ff_ram[6603] = 8'h20;
    ff_ram[6604] = 8'h20;
    ff_ram[6605] = 8'h20;
    ff_ram[6606] = 8'h20;
    ff_ram[6607] = 8'h20;
    ff_ram[6608] = 8'h20;
    ff_ram[6609] = 8'h20;
    ff_ram[6610] = 8'h20;
    ff_ram[6611] = 8'h20;
    ff_ram[6612] = 8'h20;
    ff_ram[6613] = 8'h20;
    ff_ram[6614] = 8'h20;
    ff_ram[6615] = 8'h20;
    ff_ram[6616] = 8'h20;
    ff_ram[6617] = 8'h20;
    ff_ram[6618] = 8'h20;
    ff_ram[6619] = 8'h20;
    ff_ram[6620] = 8'h20;
    ff_ram[6621] = 8'h20;
    ff_ram[6622] = 8'h20;
    ff_ram[6623] = 8'h20;
    ff_ram[6624] = 8'h20;
    ff_ram[6625] = 8'h20;
    ff_ram[6626] = 8'h20;
    ff_ram[6627] = 8'h20;
    ff_ram[6628] = 8'h20;
    ff_ram[6629] = 8'h20;
    ff_ram[6630] = 8'h20;
    ff_ram[6631] = 8'h20;
    ff_ram[6632] = 8'h20;
    ff_ram[6633] = 8'h20;
    ff_ram[6634] = 8'h20;
    ff_ram[6635] = 8'h20;
    ff_ram[6636] = 8'h20;
    ff_ram[6637] = 8'h20;
    ff_ram[6638] = 8'h20;
    ff_ram[6639] = 8'h20;
    ff_ram[6640] = 8'h20;
    ff_ram[6641] = 8'h20;
    ff_ram[6642] = 8'h20;
    ff_ram[6643] = 8'h20;
    ff_ram[6644] = 8'h20;
    ff_ram[6645] = 8'h20;
    ff_ram[6646] = 8'h20;
    ff_ram[6647] = 8'h20;
    ff_ram[6648] = 8'h20;
    ff_ram[6649] = 8'h20;
    ff_ram[6650] = 8'h20;
    ff_ram[6651] = 8'h20;
    ff_ram[6652] = 8'h20;
    ff_ram[6653] = 8'h20;
    ff_ram[6654] = 8'h20;
    ff_ram[6655] = 8'h20;
    ff_ram[6656] = 8'h20;
    ff_ram[6657] = 8'h20;
    ff_ram[6658] = 8'h20;
    ff_ram[6659] = 8'h20;
    ff_ram[6660] = 8'h20;
    ff_ram[6661] = 8'h20;
    ff_ram[6662] = 8'h20;
    ff_ram[6663] = 8'h20;
    ff_ram[6664] = 8'h20;
    ff_ram[6665] = 8'h20;
    ff_ram[6666] = 8'h20;
    ff_ram[6667] = 8'h20;
    ff_ram[6668] = 8'h20;
    ff_ram[6669] = 8'h20;
    ff_ram[6670] = 8'h20;
    ff_ram[6671] = 8'h20;
    ff_ram[6672] = 8'h20;
    ff_ram[6673] = 8'h20;
    ff_ram[6674] = 8'h20;
    ff_ram[6675] = 8'h20;
    ff_ram[6676] = 8'h20;
    ff_ram[6677] = 8'h20;
    ff_ram[6678] = 8'h20;
    ff_ram[6679] = 8'h20;
    ff_ram[6680] = 8'h20;
    ff_ram[6681] = 8'h20;
    ff_ram[6682] = 8'h20;
    ff_ram[6683] = 8'h20;
    ff_ram[6684] = 8'h20;
    ff_ram[6685] = 8'h20;
    ff_ram[6686] = 8'h20;
    ff_ram[6687] = 8'h20;
    ff_ram[6688] = 8'h20;
    ff_ram[6689] = 8'h20;
    ff_ram[6690] = 8'h20;
    ff_ram[6691] = 8'h20;
    ff_ram[6692] = 8'h20;
    ff_ram[6693] = 8'h20;
    ff_ram[6694] = 8'h20;
    ff_ram[6695] = 8'h20;
    ff_ram[6696] = 8'h20;
    ff_ram[6697] = 8'h20;
    ff_ram[6698] = 8'h20;
    ff_ram[6699] = 8'h20;
    ff_ram[6700] = 8'h20;
    ff_ram[6701] = 8'h20;
    ff_ram[6702] = 8'h20;
    ff_ram[6703] = 8'h20;
    ff_ram[6704] = 8'h20;
    ff_ram[6705] = 8'h20;
    ff_ram[6706] = 8'h20;
    ff_ram[6707] = 8'h20;
    ff_ram[6708] = 8'h20;
    ff_ram[6709] = 8'h20;
    ff_ram[6710] = 8'h20;
    ff_ram[6711] = 8'h20;
    ff_ram[6712] = 8'h20;
    ff_ram[6713] = 8'h20;
    ff_ram[6714] = 8'h20;
    ff_ram[6715] = 8'h20;
    ff_ram[6716] = 8'h20;
    ff_ram[6717] = 8'h20;
    ff_ram[6718] = 8'h20;
    ff_ram[6719] = 8'h20;
    ff_ram[6720] = 8'h20;
    ff_ram[6721] = 8'h20;
    ff_ram[6722] = 8'h20;
    ff_ram[6723] = 8'h20;
    ff_ram[6724] = 8'h20;
    ff_ram[6725] = 8'h20;
    ff_ram[6726] = 8'h20;
    ff_ram[6727] = 8'h20;
    ff_ram[6728] = 8'h20;
    ff_ram[6729] = 8'h20;
    ff_ram[6730] = 8'h20;
    ff_ram[6731] = 8'h20;
    ff_ram[6732] = 8'h20;
    ff_ram[6733] = 8'h20;
    ff_ram[6734] = 8'h20;
    ff_ram[6735] = 8'h20;
    ff_ram[6736] = 8'h20;
    ff_ram[6737] = 8'h20;
    ff_ram[6738] = 8'h20;
    ff_ram[6739] = 8'h20;
    ff_ram[6740] = 8'h20;
    ff_ram[6741] = 8'h20;
    ff_ram[6742] = 8'h20;
    ff_ram[6743] = 8'h20;
    ff_ram[6744] = 8'h20;
    ff_ram[6745] = 8'h20;
    ff_ram[6746] = 8'h20;
    ff_ram[6747] = 8'h20;
    ff_ram[6748] = 8'h20;
    ff_ram[6749] = 8'h20;
    ff_ram[6750] = 8'h20;
    ff_ram[6751] = 8'h20;
    ff_ram[6752] = 8'h20;
    ff_ram[6753] = 8'h20;
    ff_ram[6754] = 8'h20;
    ff_ram[6755] = 8'h20;
    ff_ram[6756] = 8'h20;
    ff_ram[6757] = 8'h20;
    ff_ram[6758] = 8'h20;
    ff_ram[6759] = 8'h20;
    ff_ram[6760] = 8'h20;
    ff_ram[6761] = 8'h20;
    ff_ram[6762] = 8'h20;
    ff_ram[6763] = 8'h20;
    ff_ram[6764] = 8'h20;
    ff_ram[6765] = 8'h20;
    ff_ram[6766] = 8'h20;
    ff_ram[6767] = 8'h20;
    ff_ram[6768] = 8'h20;
    ff_ram[6769] = 8'h20;
    ff_ram[6770] = 8'h20;
    ff_ram[6771] = 8'h20;
    ff_ram[6772] = 8'h20;
    ff_ram[6773] = 8'h20;
    ff_ram[6774] = 8'h20;
    ff_ram[6775] = 8'h20;
    ff_ram[6776] = 8'h20;
    ff_ram[6777] = 8'h20;
    ff_ram[6778] = 8'h20;
    ff_ram[6779] = 8'h20;
    ff_ram[6780] = 8'h20;
    ff_ram[6781] = 8'h20;
    ff_ram[6782] = 8'h20;
    ff_ram[6783] = 8'h20;
    ff_ram[6784] = 8'h20;
    ff_ram[6785] = 8'h20;
    ff_ram[6786] = 8'h20;
    ff_ram[6787] = 8'h20;
    ff_ram[6788] = 8'h20;
    ff_ram[6789] = 8'h20;
    ff_ram[6790] = 8'h20;
    ff_ram[6791] = 8'h20;
    ff_ram[6792] = 8'h20;
    ff_ram[6793] = 8'h20;
    ff_ram[6794] = 8'h20;
    ff_ram[6795] = 8'h20;
    ff_ram[6796] = 8'h20;
    ff_ram[6797] = 8'h20;
    ff_ram[6798] = 8'h20;
    ff_ram[6799] = 8'h20;
    ff_ram[6800] = 8'h20;
    ff_ram[6801] = 8'h20;
    ff_ram[6802] = 8'h20;
    ff_ram[6803] = 8'h20;
    ff_ram[6804] = 8'h20;
    ff_ram[6805] = 8'h20;
    ff_ram[6806] = 8'h20;
    ff_ram[6807] = 8'h20;
    ff_ram[6808] = 8'h20;
    ff_ram[6809] = 8'h20;
    ff_ram[6810] = 8'h20;
    ff_ram[6811] = 8'h20;
    ff_ram[6812] = 8'h20;
    ff_ram[6813] = 8'h20;
    ff_ram[6814] = 8'h20;
    ff_ram[6815] = 8'h20;
    ff_ram[6816] = 8'h20;
    ff_ram[6817] = 8'h20;
    ff_ram[6818] = 8'h20;
    ff_ram[6819] = 8'h20;
    ff_ram[6820] = 8'h20;
    ff_ram[6821] = 8'h20;
    ff_ram[6822] = 8'h20;
    ff_ram[6823] = 8'h20;
    ff_ram[6824] = 8'h20;
    ff_ram[6825] = 8'h20;
    ff_ram[6826] = 8'h20;
    ff_ram[6827] = 8'h20;
    ff_ram[6828] = 8'h20;
    ff_ram[6829] = 8'h20;
    ff_ram[6830] = 8'h20;
    ff_ram[6831] = 8'h20;
    ff_ram[6832] = 8'h20;
    ff_ram[6833] = 8'h20;
    ff_ram[6834] = 8'h20;
    ff_ram[6835] = 8'h20;
    ff_ram[6836] = 8'h20;
    ff_ram[6837] = 8'h20;
    ff_ram[6838] = 8'h20;
    ff_ram[6839] = 8'h20;
    ff_ram[6840] = 8'h20;
    ff_ram[6841] = 8'h20;
    ff_ram[6842] = 8'h20;
    ff_ram[6843] = 8'h20;
    ff_ram[6844] = 8'h20;
    ff_ram[6845] = 8'h20;
    ff_ram[6846] = 8'h20;
    ff_ram[6847] = 8'h20;
    ff_ram[6848] = 8'h20;
    ff_ram[6849] = 8'h20;
    ff_ram[6850] = 8'h20;
    ff_ram[6851] = 8'h20;
    ff_ram[6852] = 8'h20;
    ff_ram[6853] = 8'h20;
    ff_ram[6854] = 8'h20;
    ff_ram[6855] = 8'h20;
    ff_ram[6856] = 8'h20;
    ff_ram[6857] = 8'h20;
    ff_ram[6858] = 8'h20;
    ff_ram[6859] = 8'h20;
    ff_ram[6860] = 8'h20;
    ff_ram[6861] = 8'h20;
    ff_ram[6862] = 8'h20;
    ff_ram[6863] = 8'h20;
    ff_ram[6864] = 8'h20;
    ff_ram[6865] = 8'h20;
    ff_ram[6866] = 8'h20;
    ff_ram[6867] = 8'h20;
    ff_ram[6868] = 8'h20;
    ff_ram[6869] = 8'h20;
    ff_ram[6870] = 8'h20;
    ff_ram[6871] = 8'h20;
    ff_ram[6872] = 8'h20;
    ff_ram[6873] = 8'h20;
    ff_ram[6874] = 8'h20;
    ff_ram[6875] = 8'h20;
    ff_ram[6876] = 8'h20;
    ff_ram[6877] = 8'h20;
    ff_ram[6878] = 8'h20;
    ff_ram[6879] = 8'h20;
    ff_ram[6880] = 8'h20;
    ff_ram[6881] = 8'h20;
    ff_ram[6882] = 8'h63;
    ff_ram[6883] = 8'h6F;
    ff_ram[6884] = 8'h6C;
    ff_ram[6885] = 8'h6F;
    ff_ram[6886] = 8'h72;
    ff_ram[6887] = 8'h20;
    ff_ram[6888] = 8'h61;
    ff_ram[6889] = 8'h75;
    ff_ram[6890] = 8'h74;
    ff_ram[6891] = 8'h6F;
    ff_ram[6892] = 8'h20;
    ff_ram[6893] = 8'h20;
    ff_ram[6894] = 8'h67;
    ff_ram[6895] = 8'h6F;
    ff_ram[6896] = 8'h74;
    ff_ram[6897] = 8'h6F;
    ff_ram[6898] = 8'h20;
    ff_ram[6899] = 8'h20;
    ff_ram[6900] = 8'h6C;
    ff_ram[6901] = 8'h69;
    ff_ram[6902] = 8'h73;
    ff_ram[6903] = 8'h74;
    ff_ram[6904] = 8'h20;
    ff_ram[6905] = 8'h20;
    ff_ram[6906] = 8'h72;
    ff_ram[6907] = 8'h75;
    ff_ram[6908] = 8'h6E;
    ff_ram[6909] = 8'h20;
    ff_ram[6910] = 8'h20;
    ff_ram[6911] = 8'h20;
    ff_ram[6912] = 8'hD1;
    ff_ram[6913] = 8'h00;
    ff_ram[6914] = 8'h00;
    ff_ram[6915] = 8'h0F;
    ff_ram[6916] = 8'hD1;
    ff_ram[6917] = 8'h00;
    ff_ram[6918] = 8'h01;
    ff_ram[6919] = 8'h0F;
    ff_ram[6920] = 8'hD1;
    ff_ram[6921] = 8'h00;
    ff_ram[6922] = 8'h02;
    ff_ram[6923] = 8'h0F;
    ff_ram[6924] = 8'hD1;
    ff_ram[6925] = 8'h00;
    ff_ram[6926] = 8'h03;
    ff_ram[6927] = 8'h0F;
    ff_ram[6928] = 8'hD1;
    ff_ram[6929] = 8'h00;
    ff_ram[6930] = 8'h04;
    ff_ram[6931] = 8'h0F;
    ff_ram[6932] = 8'hD1;
    ff_ram[6933] = 8'h00;
    ff_ram[6934] = 8'h05;
    ff_ram[6935] = 8'h0F;
    ff_ram[6936] = 8'hD1;
    ff_ram[6937] = 8'h00;
    ff_ram[6938] = 8'h06;
    ff_ram[6939] = 8'h0F;
    ff_ram[6940] = 8'hD1;
    ff_ram[6941] = 8'h00;
    ff_ram[6942] = 8'h07;
    ff_ram[6943] = 8'h0F;
    ff_ram[6944] = 8'hD1;
    ff_ram[6945] = 8'h00;
    ff_ram[6946] = 8'h08;
    ff_ram[6947] = 8'h0F;
    ff_ram[6948] = 8'hD1;
    ff_ram[6949] = 8'h00;
    ff_ram[6950] = 8'h09;
    ff_ram[6951] = 8'h0F;
    ff_ram[6952] = 8'hD1;
    ff_ram[6953] = 8'h00;
    ff_ram[6954] = 8'h0A;
    ff_ram[6955] = 8'h0F;
    ff_ram[6956] = 8'hD1;
    ff_ram[6957] = 8'h00;
    ff_ram[6958] = 8'h0B;
    ff_ram[6959] = 8'h0F;
    ff_ram[6960] = 8'hD1;
    ff_ram[6961] = 8'h00;
    ff_ram[6962] = 8'h0C;
    ff_ram[6963] = 8'h0F;
    ff_ram[6964] = 8'hD1;
    ff_ram[6965] = 8'h00;
    ff_ram[6966] = 8'h0D;
    ff_ram[6967] = 8'h0F;
    ff_ram[6968] = 8'hD1;
    ff_ram[6969] = 8'h00;
    ff_ram[6970] = 8'h0E;
    ff_ram[6971] = 8'h0F;
    ff_ram[6972] = 8'hD1;
    ff_ram[6973] = 8'h00;
    ff_ram[6974] = 8'h0F;
    ff_ram[6975] = 8'h0F;
    ff_ram[6976] = 8'hD1;
    ff_ram[6977] = 8'h00;
    ff_ram[6978] = 8'h10;
    ff_ram[6979] = 8'h0F;
    ff_ram[6980] = 8'hD1;
    ff_ram[6981] = 8'h00;
    ff_ram[6982] = 8'h11;
    ff_ram[6983] = 8'h0F;
    ff_ram[6984] = 8'hD1;
    ff_ram[6985] = 8'h00;
    ff_ram[6986] = 8'h12;
    ff_ram[6987] = 8'h0F;
    ff_ram[6988] = 8'hD1;
    ff_ram[6989] = 8'h00;
    ff_ram[6990] = 8'h13;
    ff_ram[6991] = 8'h0F;
    ff_ram[6992] = 8'hD1;
    ff_ram[6993] = 8'h00;
    ff_ram[6994] = 8'h14;
    ff_ram[6995] = 8'h0F;
    ff_ram[6996] = 8'hD1;
    ff_ram[6997] = 8'h00;
    ff_ram[6998] = 8'h15;
    ff_ram[6999] = 8'h0F;
    ff_ram[7000] = 8'hD1;
    ff_ram[7001] = 8'h00;
    ff_ram[7002] = 8'h16;
    ff_ram[7003] = 8'h0F;
    ff_ram[7004] = 8'hD1;
    ff_ram[7005] = 8'h00;
    ff_ram[7006] = 8'h17;
    ff_ram[7007] = 8'h0F;
    ff_ram[7008] = 8'hD1;
    ff_ram[7009] = 8'h00;
    ff_ram[7010] = 8'h18;
    ff_ram[7011] = 8'h0F;
    ff_ram[7012] = 8'hD1;
    ff_ram[7013] = 8'h00;
    ff_ram[7014] = 8'h19;
    ff_ram[7015] = 8'h0F;
    ff_ram[7016] = 8'hD1;
    ff_ram[7017] = 8'h00;
    ff_ram[7018] = 8'h1A;
    ff_ram[7019] = 8'h0F;
    ff_ram[7020] = 8'hD1;
    ff_ram[7021] = 8'h00;
    ff_ram[7022] = 8'h1B;
    ff_ram[7023] = 8'h0F;
    ff_ram[7024] = 8'hD1;
    ff_ram[7025] = 8'h00;
    ff_ram[7026] = 8'h1C;
    ff_ram[7027] = 8'h0F;
    ff_ram[7028] = 8'hD1;
    ff_ram[7029] = 8'h00;
    ff_ram[7030] = 8'h1D;
    ff_ram[7031] = 8'h0F;
    ff_ram[7032] = 8'hD1;
    ff_ram[7033] = 8'h00;
    ff_ram[7034] = 8'h1E;
    ff_ram[7035] = 8'h0F;
    ff_ram[7036] = 8'hD1;
    ff_ram[7037] = 8'h00;
    ff_ram[7038] = 8'h1F;
    ff_ram[7039] = 8'h0F;
    ff_ram[7040] = 8'h00;
    ff_ram[7041] = 8'h00;
    ff_ram[7042] = 8'h00;
    ff_ram[7043] = 8'h00;
    ff_ram[7044] = 8'h11;
    ff_ram[7045] = 8'h06;
    ff_ram[7046] = 8'h33;
    ff_ram[7047] = 8'h07;
    ff_ram[7048] = 8'h17;
    ff_ram[7049] = 8'h01;
    ff_ram[7050] = 8'h27;
    ff_ram[7051] = 8'h03;
    ff_ram[7052] = 8'h51;
    ff_ram[7053] = 8'h01;
    ff_ram[7054] = 8'h27;
    ff_ram[7055] = 8'h06;
    ff_ram[7056] = 8'h71;
    ff_ram[7057] = 8'h01;
    ff_ram[7058] = 8'h73;
    ff_ram[7059] = 8'h03;
    ff_ram[7060] = 8'h61;
    ff_ram[7061] = 8'h06;
    ff_ram[7062] = 8'h64;
    ff_ram[7063] = 8'h06;
    ff_ram[7064] = 8'h11;
    ff_ram[7065] = 8'h04;
    ff_ram[7066] = 8'h65;
    ff_ram[7067] = 8'h02;
    ff_ram[7068] = 8'h55;
    ff_ram[7069] = 8'h05;
    ff_ram[7070] = 8'h77;
    ff_ram[7071] = 8'h07;
    ff_ram[7072] = 8'h00;
    ff_ram[7073] = 8'h00;
    ff_ram[7074] = 8'h00;
    ff_ram[7075] = 8'h00;
    ff_ram[7076] = 8'h00;
    ff_ram[7077] = 8'h00;
    ff_ram[7078] = 8'h00;
    ff_ram[7079] = 8'h00;
    ff_ram[7080] = 8'h00;
    ff_ram[7081] = 8'h00;
    ff_ram[7082] = 8'h00;
    ff_ram[7083] = 8'h00;
    ff_ram[7084] = 8'h00;
    ff_ram[7085] = 8'h00;
    ff_ram[7086] = 8'h00;
    ff_ram[7087] = 8'h00;
    ff_ram[7088] = 8'h00;
    ff_ram[7089] = 8'h00;
    ff_ram[7090] = 8'h00;
    ff_ram[7091] = 8'h00;
    ff_ram[7092] = 8'h00;
    ff_ram[7093] = 8'h00;
    ff_ram[7094] = 8'h00;
    ff_ram[7095] = 8'h00;
    ff_ram[7096] = 8'h00;
    ff_ram[7097] = 8'h00;
    ff_ram[7098] = 8'h00;
    ff_ram[7099] = 8'h00;
    ff_ram[7100] = 8'h00;
    ff_ram[7101] = 8'h00;
    ff_ram[7102] = 8'h00;
    ff_ram[7103] = 8'h00;
    ff_ram[7104] = 8'h00;
    ff_ram[7105] = 8'h00;
    ff_ram[7106] = 8'h00;
    ff_ram[7107] = 8'h00;
    ff_ram[7108] = 8'h00;
    ff_ram[7109] = 8'h00;
    ff_ram[7110] = 8'h00;
    ff_ram[7111] = 8'h00;
    ff_ram[7112] = 8'h00;
    ff_ram[7113] = 8'h00;
    ff_ram[7114] = 8'h00;
    ff_ram[7115] = 8'h00;
    ff_ram[7116] = 8'h00;
    ff_ram[7117] = 8'h00;
    ff_ram[7118] = 8'h00;
    ff_ram[7119] = 8'h00;
    ff_ram[7120] = 8'h00;
    ff_ram[7121] = 8'h00;
    ff_ram[7122] = 8'h00;
    ff_ram[7123] = 8'h00;
    ff_ram[7124] = 8'h00;
    ff_ram[7125] = 8'h00;
    ff_ram[7126] = 8'h00;
    ff_ram[7127] = 8'h00;
    ff_ram[7128] = 8'h00;
    ff_ram[7129] = 8'h00;
    ff_ram[7130] = 8'h00;
    ff_ram[7131] = 8'h00;
    ff_ram[7132] = 8'h00;
    ff_ram[7133] = 8'h00;
    ff_ram[7134] = 8'h00;
    ff_ram[7135] = 8'h00;
    ff_ram[7136] = 8'h00;
    ff_ram[7137] = 8'h00;
    ff_ram[7138] = 8'h00;
    ff_ram[7139] = 8'h00;
    ff_ram[7140] = 8'h00;
    ff_ram[7141] = 8'h00;
    ff_ram[7142] = 8'h00;
    ff_ram[7143] = 8'h00;
    ff_ram[7144] = 8'h00;
    ff_ram[7145] = 8'h00;
    ff_ram[7146] = 8'h00;
    ff_ram[7147] = 8'h00;
    ff_ram[7148] = 8'h00;
    ff_ram[7149] = 8'h00;
    ff_ram[7150] = 8'h00;
    ff_ram[7151] = 8'h00;
    ff_ram[7152] = 8'h00;
    ff_ram[7153] = 8'h00;
    ff_ram[7154] = 8'h00;
    ff_ram[7155] = 8'h00;
    ff_ram[7156] = 8'h00;
    ff_ram[7157] = 8'h00;
    ff_ram[7158] = 8'h00;
    ff_ram[7159] = 8'h00;
    ff_ram[7160] = 8'h00;
    ff_ram[7161] = 8'h00;
    ff_ram[7162] = 8'h00;
    ff_ram[7163] = 8'h00;
    ff_ram[7164] = 8'h00;
    ff_ram[7165] = 8'h00;
    ff_ram[7166] = 8'h00;
    ff_ram[7167] = 8'h00;
    ff_ram[7168] = 8'h00;
    ff_ram[7169] = 8'h00;
    ff_ram[7170] = 8'h00;
    ff_ram[7171] = 8'h00;
    ff_ram[7172] = 8'h00;
    ff_ram[7173] = 8'h00;
    ff_ram[7174] = 8'h00;
    ff_ram[7175] = 8'h00;
    ff_ram[7176] = 8'h00;
    ff_ram[7177] = 8'h00;
    ff_ram[7178] = 8'h00;
    ff_ram[7179] = 8'h00;
    ff_ram[7180] = 8'h00;
    ff_ram[7181] = 8'h00;
    ff_ram[7182] = 8'h00;
    ff_ram[7183] = 8'h00;
    ff_ram[7184] = 8'h00;
    ff_ram[7185] = 8'h00;
    ff_ram[7186] = 8'h00;
    ff_ram[7187] = 8'h00;
    ff_ram[7188] = 8'h00;
    ff_ram[7189] = 8'h00;
    ff_ram[7190] = 8'h00;
    ff_ram[7191] = 8'h00;
    ff_ram[7192] = 8'h00;
    ff_ram[7193] = 8'h00;
    ff_ram[7194] = 8'h00;
    ff_ram[7195] = 8'h00;
    ff_ram[7196] = 8'h00;
    ff_ram[7197] = 8'h00;
    ff_ram[7198] = 8'h00;
    ff_ram[7199] = 8'h00;
    ff_ram[7200] = 8'h00;
    ff_ram[7201] = 8'h00;
    ff_ram[7202] = 8'h00;
    ff_ram[7203] = 8'h00;
    ff_ram[7204] = 8'h00;
    ff_ram[7205] = 8'h00;
    ff_ram[7206] = 8'h00;
    ff_ram[7207] = 8'h00;
    ff_ram[7208] = 8'h00;
    ff_ram[7209] = 8'h00;
    ff_ram[7210] = 8'h00;
    ff_ram[7211] = 8'h00;
    ff_ram[7212] = 8'h00;
    ff_ram[7213] = 8'h00;
    ff_ram[7214] = 8'h00;
    ff_ram[7215] = 8'h00;
    ff_ram[7216] = 8'h00;
    ff_ram[7217] = 8'h00;
    ff_ram[7218] = 8'h00;
    ff_ram[7219] = 8'h00;
    ff_ram[7220] = 8'h00;
    ff_ram[7221] = 8'h00;
    ff_ram[7222] = 8'h00;
    ff_ram[7223] = 8'h00;
    ff_ram[7224] = 8'h00;
    ff_ram[7225] = 8'h00;
    ff_ram[7226] = 8'h00;
    ff_ram[7227] = 8'h00;
    ff_ram[7228] = 8'h00;
    ff_ram[7229] = 8'h00;
    ff_ram[7230] = 8'h00;
    ff_ram[7231] = 8'h00;
    ff_ram[7232] = 8'h00;
    ff_ram[7233] = 8'h00;
    ff_ram[7234] = 8'h00;
    ff_ram[7235] = 8'h00;
    ff_ram[7236] = 8'h00;
    ff_ram[7237] = 8'h00;
    ff_ram[7238] = 8'h00;
    ff_ram[7239] = 8'h00;
    ff_ram[7240] = 8'h00;
    ff_ram[7241] = 8'h00;
    ff_ram[7242] = 8'h00;
    ff_ram[7243] = 8'h00;
    ff_ram[7244] = 8'h00;
    ff_ram[7245] = 8'h00;
    ff_ram[7246] = 8'h00;
    ff_ram[7247] = 8'h00;
    ff_ram[7248] = 8'h00;
    ff_ram[7249] = 8'h00;
    ff_ram[7250] = 8'h00;
    ff_ram[7251] = 8'h00;
    ff_ram[7252] = 8'h00;
    ff_ram[7253] = 8'h00;
    ff_ram[7254] = 8'h00;
    ff_ram[7255] = 8'h00;
    ff_ram[7256] = 8'h00;
    ff_ram[7257] = 8'h00;
    ff_ram[7258] = 8'h00;
    ff_ram[7259] = 8'h00;
    ff_ram[7260] = 8'h00;
    ff_ram[7261] = 8'h00;
    ff_ram[7262] = 8'h00;
    ff_ram[7263] = 8'h00;
    ff_ram[7264] = 8'h00;
    ff_ram[7265] = 8'h00;
    ff_ram[7266] = 8'h00;
    ff_ram[7267] = 8'h00;
    ff_ram[7268] = 8'h00;
    ff_ram[7269] = 8'h00;
    ff_ram[7270] = 8'h00;
    ff_ram[7271] = 8'h00;
    ff_ram[7272] = 8'h00;
    ff_ram[7273] = 8'h00;
    ff_ram[7274] = 8'h00;
    ff_ram[7275] = 8'h00;
    ff_ram[7276] = 8'h00;
    ff_ram[7277] = 8'h00;
    ff_ram[7278] = 8'h00;
    ff_ram[7279] = 8'h00;
    ff_ram[7280] = 8'h00;
    ff_ram[7281] = 8'h00;
    ff_ram[7282] = 8'h00;
    ff_ram[7283] = 8'h00;
    ff_ram[7284] = 8'h00;
    ff_ram[7285] = 8'h00;
    ff_ram[7286] = 8'h00;
    ff_ram[7287] = 8'h00;
    ff_ram[7288] = 8'h00;
    ff_ram[7289] = 8'h00;
    ff_ram[7290] = 8'h00;
    ff_ram[7291] = 8'h00;
    ff_ram[7292] = 8'h00;
    ff_ram[7293] = 8'h00;
    ff_ram[7294] = 8'h00;
    ff_ram[7295] = 8'h00;
    ff_ram[7296] = 8'h00;
    ff_ram[7297] = 8'h00;
    ff_ram[7298] = 8'h00;
    ff_ram[7299] = 8'h00;
    ff_ram[7300] = 8'h00;
    ff_ram[7301] = 8'h00;
    ff_ram[7302] = 8'h00;
    ff_ram[7303] = 8'h00;
    ff_ram[7304] = 8'h00;
    ff_ram[7305] = 8'h00;
    ff_ram[7306] = 8'h00;
    ff_ram[7307] = 8'h00;
    ff_ram[7308] = 8'h00;
    ff_ram[7309] = 8'h00;
    ff_ram[7310] = 8'h00;
    ff_ram[7311] = 8'h00;
    ff_ram[7312] = 8'h00;
    ff_ram[7313] = 8'h00;
    ff_ram[7314] = 8'h00;
    ff_ram[7315] = 8'h00;
    ff_ram[7316] = 8'h00;
    ff_ram[7317] = 8'h00;
    ff_ram[7318] = 8'h00;
    ff_ram[7319] = 8'h00;
    ff_ram[7320] = 8'h00;
    ff_ram[7321] = 8'h00;
    ff_ram[7322] = 8'h00;
    ff_ram[7323] = 8'h00;
    ff_ram[7324] = 8'h00;
    ff_ram[7325] = 8'h00;
    ff_ram[7326] = 8'h00;
    ff_ram[7327] = 8'h00;
    ff_ram[7328] = 8'h00;
    ff_ram[7329] = 8'h00;
    ff_ram[7330] = 8'h00;
    ff_ram[7331] = 8'h00;
    ff_ram[7332] = 8'h00;
    ff_ram[7333] = 8'h00;
    ff_ram[7334] = 8'h00;
    ff_ram[7335] = 8'h00;
    ff_ram[7336] = 8'h00;
    ff_ram[7337] = 8'h00;
    ff_ram[7338] = 8'h00;
    ff_ram[7339] = 8'h00;
    ff_ram[7340] = 8'h00;
    ff_ram[7341] = 8'h00;
    ff_ram[7342] = 8'h00;
    ff_ram[7343] = 8'h00;
    ff_ram[7344] = 8'h00;
    ff_ram[7345] = 8'h00;
    ff_ram[7346] = 8'h00;
    ff_ram[7347] = 8'h00;
    ff_ram[7348] = 8'h00;
    ff_ram[7349] = 8'h00;
    ff_ram[7350] = 8'h00;
    ff_ram[7351] = 8'h00;
    ff_ram[7352] = 8'h00;
    ff_ram[7353] = 8'h00;
    ff_ram[7354] = 8'h00;
    ff_ram[7355] = 8'h00;
    ff_ram[7356] = 8'h00;
    ff_ram[7357] = 8'h00;
    ff_ram[7358] = 8'h00;
    ff_ram[7359] = 8'h00;
    ff_ram[7360] = 8'h00;
    ff_ram[7361] = 8'h00;
    ff_ram[7362] = 8'h00;
    ff_ram[7363] = 8'h00;
    ff_ram[7364] = 8'h00;
    ff_ram[7365] = 8'h00;
    ff_ram[7366] = 8'h00;
    ff_ram[7367] = 8'h00;
    ff_ram[7368] = 8'h00;
    ff_ram[7369] = 8'h00;
    ff_ram[7370] = 8'h00;
    ff_ram[7371] = 8'h00;
    ff_ram[7372] = 8'h00;
    ff_ram[7373] = 8'h00;
    ff_ram[7374] = 8'h00;
    ff_ram[7375] = 8'h00;
    ff_ram[7376] = 8'h00;
    ff_ram[7377] = 8'h00;
    ff_ram[7378] = 8'h00;
    ff_ram[7379] = 8'h00;
    ff_ram[7380] = 8'h00;
    ff_ram[7381] = 8'h00;
    ff_ram[7382] = 8'h00;
    ff_ram[7383] = 8'h00;
    ff_ram[7384] = 8'h00;
    ff_ram[7385] = 8'h00;
    ff_ram[7386] = 8'h00;
    ff_ram[7387] = 8'h00;
    ff_ram[7388] = 8'h00;
    ff_ram[7389] = 8'h00;
    ff_ram[7390] = 8'h00;
    ff_ram[7391] = 8'h00;
    ff_ram[7392] = 8'h00;
    ff_ram[7393] = 8'h00;
    ff_ram[7394] = 8'h00;
    ff_ram[7395] = 8'h00;
    ff_ram[7396] = 8'h00;
    ff_ram[7397] = 8'h00;
    ff_ram[7398] = 8'h00;
    ff_ram[7399] = 8'h00;
    ff_ram[7400] = 8'h00;
    ff_ram[7401] = 8'h00;
    ff_ram[7402] = 8'h00;
    ff_ram[7403] = 8'h00;
    ff_ram[7404] = 8'h00;
    ff_ram[7405] = 8'h00;
    ff_ram[7406] = 8'h00;
    ff_ram[7407] = 8'h00;
    ff_ram[7408] = 8'h00;
    ff_ram[7409] = 8'h00;
    ff_ram[7410] = 8'h00;
    ff_ram[7411] = 8'h00;
    ff_ram[7412] = 8'h00;
    ff_ram[7413] = 8'h00;
    ff_ram[7414] = 8'h00;
    ff_ram[7415] = 8'h00;
    ff_ram[7416] = 8'h00;
    ff_ram[7417] = 8'h00;
    ff_ram[7418] = 8'h00;
    ff_ram[7419] = 8'h00;
    ff_ram[7420] = 8'h00;
    ff_ram[7421] = 8'h00;
    ff_ram[7422] = 8'h00;
    ff_ram[7423] = 8'h00;
    ff_ram[7424] = 8'h00;
    ff_ram[7425] = 8'h00;
    ff_ram[7426] = 8'h00;
    ff_ram[7427] = 8'h00;
    ff_ram[7428] = 8'h00;
    ff_ram[7429] = 8'h00;
    ff_ram[7430] = 8'h00;
    ff_ram[7431] = 8'h00;
    ff_ram[7432] = 8'h00;
    ff_ram[7433] = 8'h00;
    ff_ram[7434] = 8'h00;
    ff_ram[7435] = 8'h00;
    ff_ram[7436] = 8'h00;
    ff_ram[7437] = 8'h00;
    ff_ram[7438] = 8'h00;
    ff_ram[7439] = 8'h00;
    ff_ram[7440] = 8'h00;
    ff_ram[7441] = 8'h00;
    ff_ram[7442] = 8'h00;
    ff_ram[7443] = 8'h00;
    ff_ram[7444] = 8'h00;
    ff_ram[7445] = 8'h00;
    ff_ram[7446] = 8'h00;
    ff_ram[7447] = 8'h00;
    ff_ram[7448] = 8'h00;
    ff_ram[7449] = 8'h00;
    ff_ram[7450] = 8'h00;
    ff_ram[7451] = 8'h00;
    ff_ram[7452] = 8'h00;
    ff_ram[7453] = 8'h00;
    ff_ram[7454] = 8'h00;
    ff_ram[7455] = 8'h00;
    ff_ram[7456] = 8'h00;
    ff_ram[7457] = 8'h00;
    ff_ram[7458] = 8'h00;
    ff_ram[7459] = 8'h00;
    ff_ram[7460] = 8'h00;
    ff_ram[7461] = 8'h00;
    ff_ram[7462] = 8'h00;
    ff_ram[7463] = 8'h00;
    ff_ram[7464] = 8'h00;
    ff_ram[7465] = 8'h00;
    ff_ram[7466] = 8'h00;
    ff_ram[7467] = 8'h00;
    ff_ram[7468] = 8'h00;
    ff_ram[7469] = 8'h00;
    ff_ram[7470] = 8'h00;
    ff_ram[7471] = 8'h00;
    ff_ram[7472] = 8'h00;
    ff_ram[7473] = 8'h00;
    ff_ram[7474] = 8'h00;
    ff_ram[7475] = 8'h00;
    ff_ram[7476] = 8'h00;
    ff_ram[7477] = 8'h00;
    ff_ram[7478] = 8'h00;
    ff_ram[7479] = 8'h00;
    ff_ram[7480] = 8'h00;
    ff_ram[7481] = 8'h00;
    ff_ram[7482] = 8'h00;
    ff_ram[7483] = 8'h00;
    ff_ram[7484] = 8'h00;
    ff_ram[7485] = 8'h00;
    ff_ram[7486] = 8'h00;
    ff_ram[7487] = 8'h00;
    ff_ram[7488] = 8'h00;
    ff_ram[7489] = 8'h00;
    ff_ram[7490] = 8'h00;
    ff_ram[7491] = 8'h00;
    ff_ram[7492] = 8'h00;
    ff_ram[7493] = 8'h00;
    ff_ram[7494] = 8'h00;
    ff_ram[7495] = 8'h00;
    ff_ram[7496] = 8'h00;
    ff_ram[7497] = 8'h00;
    ff_ram[7498] = 8'h00;
    ff_ram[7499] = 8'h00;
    ff_ram[7500] = 8'h00;
    ff_ram[7501] = 8'h00;
    ff_ram[7502] = 8'h00;
    ff_ram[7503] = 8'h00;
    ff_ram[7504] = 8'h00;
    ff_ram[7505] = 8'h00;
    ff_ram[7506] = 8'h00;
    ff_ram[7507] = 8'h00;
    ff_ram[7508] = 8'h00;
    ff_ram[7509] = 8'h00;
    ff_ram[7510] = 8'h00;
    ff_ram[7511] = 8'h00;
    ff_ram[7512] = 8'h00;
    ff_ram[7513] = 8'h00;
    ff_ram[7514] = 8'h00;
    ff_ram[7515] = 8'h00;
    ff_ram[7516] = 8'h00;
    ff_ram[7517] = 8'h00;
    ff_ram[7518] = 8'h00;
    ff_ram[7519] = 8'h00;
    ff_ram[7520] = 8'h00;
    ff_ram[7521] = 8'h00;
    ff_ram[7522] = 8'h00;
    ff_ram[7523] = 8'h00;
    ff_ram[7524] = 8'h00;
    ff_ram[7525] = 8'h00;
    ff_ram[7526] = 8'h00;
    ff_ram[7527] = 8'h00;
    ff_ram[7528] = 8'h00;
    ff_ram[7529] = 8'h00;
    ff_ram[7530] = 8'h00;
    ff_ram[7531] = 8'h00;
    ff_ram[7532] = 8'h00;
    ff_ram[7533] = 8'h00;
    ff_ram[7534] = 8'h00;
    ff_ram[7535] = 8'h00;
    ff_ram[7536] = 8'h00;
    ff_ram[7537] = 8'h00;
    ff_ram[7538] = 8'h00;
    ff_ram[7539] = 8'h00;
    ff_ram[7540] = 8'h00;
    ff_ram[7541] = 8'h00;
    ff_ram[7542] = 8'h00;
    ff_ram[7543] = 8'h00;
    ff_ram[7544] = 8'h00;
    ff_ram[7545] = 8'h00;
    ff_ram[7546] = 8'h00;
    ff_ram[7547] = 8'h00;
    ff_ram[7548] = 8'h00;
    ff_ram[7549] = 8'h00;
    ff_ram[7550] = 8'h00;
    ff_ram[7551] = 8'h00;
    ff_ram[7552] = 8'h00;
    ff_ram[7553] = 8'h00;
    ff_ram[7554] = 8'h00;
    ff_ram[7555] = 8'h00;
    ff_ram[7556] = 8'h00;
    ff_ram[7557] = 8'h00;
    ff_ram[7558] = 8'h00;
    ff_ram[7559] = 8'h00;
    ff_ram[7560] = 8'h00;
    ff_ram[7561] = 8'h00;
    ff_ram[7562] = 8'h00;
    ff_ram[7563] = 8'h00;
    ff_ram[7564] = 8'h00;
    ff_ram[7565] = 8'h00;
    ff_ram[7566] = 8'h00;
    ff_ram[7567] = 8'h00;
    ff_ram[7568] = 8'h00;
    ff_ram[7569] = 8'h00;
    ff_ram[7570] = 8'h00;
    ff_ram[7571] = 8'h00;
    ff_ram[7572] = 8'h00;
    ff_ram[7573] = 8'h00;
    ff_ram[7574] = 8'h00;
    ff_ram[7575] = 8'h00;
    ff_ram[7576] = 8'h00;
    ff_ram[7577] = 8'h00;
    ff_ram[7578] = 8'h00;
    ff_ram[7579] = 8'h00;
    ff_ram[7580] = 8'h00;
    ff_ram[7581] = 8'h00;
    ff_ram[7582] = 8'h00;
    ff_ram[7583] = 8'h00;
    ff_ram[7584] = 8'h00;
    ff_ram[7585] = 8'h00;
    ff_ram[7586] = 8'h00;
    ff_ram[7587] = 8'h00;
    ff_ram[7588] = 8'h00;
    ff_ram[7589] = 8'h00;
    ff_ram[7590] = 8'h00;
    ff_ram[7591] = 8'h00;
    ff_ram[7592] = 8'h00;
    ff_ram[7593] = 8'h00;
    ff_ram[7594] = 8'h00;
    ff_ram[7595] = 8'h00;
    ff_ram[7596] = 8'h00;
    ff_ram[7597] = 8'h00;
    ff_ram[7598] = 8'h00;
    ff_ram[7599] = 8'h00;
    ff_ram[7600] = 8'h00;
    ff_ram[7601] = 8'h00;
    ff_ram[7602] = 8'h00;
    ff_ram[7603] = 8'h00;
    ff_ram[7604] = 8'h00;
    ff_ram[7605] = 8'h00;
    ff_ram[7606] = 8'h00;
    ff_ram[7607] = 8'h00;
    ff_ram[7608] = 8'h00;
    ff_ram[7609] = 8'h00;
    ff_ram[7610] = 8'h00;
    ff_ram[7611] = 8'h00;
    ff_ram[7612] = 8'h00;
    ff_ram[7613] = 8'h00;
    ff_ram[7614] = 8'h00;
    ff_ram[7615] = 8'h00;
    ff_ram[7616] = 8'h00;
    ff_ram[7617] = 8'h00;
    ff_ram[7618] = 8'h00;
    ff_ram[7619] = 8'h00;
    ff_ram[7620] = 8'h00;
    ff_ram[7621] = 8'h00;
    ff_ram[7622] = 8'h00;
    ff_ram[7623] = 8'h00;
    ff_ram[7624] = 8'h00;
    ff_ram[7625] = 8'h00;
    ff_ram[7626] = 8'h00;
    ff_ram[7627] = 8'h00;
    ff_ram[7628] = 8'h00;
    ff_ram[7629] = 8'h00;
    ff_ram[7630] = 8'h00;
    ff_ram[7631] = 8'h00;
    ff_ram[7632] = 8'h00;
    ff_ram[7633] = 8'h00;
    ff_ram[7634] = 8'h00;
    ff_ram[7635] = 8'h00;
    ff_ram[7636] = 8'h00;
    ff_ram[7637] = 8'h00;
    ff_ram[7638] = 8'h00;
    ff_ram[7639] = 8'h00;
    ff_ram[7640] = 8'h00;
    ff_ram[7641] = 8'h00;
    ff_ram[7642] = 8'h00;
    ff_ram[7643] = 8'h00;
    ff_ram[7644] = 8'h00;
    ff_ram[7645] = 8'h00;
    ff_ram[7646] = 8'h00;
    ff_ram[7647] = 8'h00;
    ff_ram[7648] = 8'h00;
    ff_ram[7649] = 8'h00;
    ff_ram[7650] = 8'h00;
    ff_ram[7651] = 8'h00;
    ff_ram[7652] = 8'h00;
    ff_ram[7653] = 8'h00;
    ff_ram[7654] = 8'h00;
    ff_ram[7655] = 8'h00;
    ff_ram[7656] = 8'h00;
    ff_ram[7657] = 8'h00;
    ff_ram[7658] = 8'h00;
    ff_ram[7659] = 8'h00;
    ff_ram[7660] = 8'h00;
    ff_ram[7661] = 8'h00;
    ff_ram[7662] = 8'h00;
    ff_ram[7663] = 8'h00;
    ff_ram[7664] = 8'h00;
    ff_ram[7665] = 8'h00;
    ff_ram[7666] = 8'h00;
    ff_ram[7667] = 8'h00;
    ff_ram[7668] = 8'h00;
    ff_ram[7669] = 8'h00;
    ff_ram[7670] = 8'h00;
    ff_ram[7671] = 8'h00;
    ff_ram[7672] = 8'h00;
    ff_ram[7673] = 8'h00;
    ff_ram[7674] = 8'h00;
    ff_ram[7675] = 8'h00;
    ff_ram[7676] = 8'h00;
    ff_ram[7677] = 8'h00;
    ff_ram[7678] = 8'h00;
    ff_ram[7679] = 8'h00;
    ff_ram[7680] = 8'h00;
    ff_ram[7681] = 8'h00;
    ff_ram[7682] = 8'h00;
    ff_ram[7683] = 8'h00;
    ff_ram[7684] = 8'h00;
    ff_ram[7685] = 8'h00;
    ff_ram[7686] = 8'h00;
    ff_ram[7687] = 8'h00;
    ff_ram[7688] = 8'h00;
    ff_ram[7689] = 8'h00;
    ff_ram[7690] = 8'h00;
    ff_ram[7691] = 8'h00;
    ff_ram[7692] = 8'h00;
    ff_ram[7693] = 8'h00;
    ff_ram[7694] = 8'h00;
    ff_ram[7695] = 8'h00;
    ff_ram[7696] = 8'h00;
    ff_ram[7697] = 8'h00;
    ff_ram[7698] = 8'h00;
    ff_ram[7699] = 8'h00;
    ff_ram[7700] = 8'h00;
    ff_ram[7701] = 8'h00;
    ff_ram[7702] = 8'h00;
    ff_ram[7703] = 8'h00;
    ff_ram[7704] = 8'h00;
    ff_ram[7705] = 8'h00;
    ff_ram[7706] = 8'h00;
    ff_ram[7707] = 8'h00;
    ff_ram[7708] = 8'h00;
    ff_ram[7709] = 8'h00;
    ff_ram[7710] = 8'h00;
    ff_ram[7711] = 8'h00;
    ff_ram[7712] = 8'h00;
    ff_ram[7713] = 8'h00;
    ff_ram[7714] = 8'h00;
    ff_ram[7715] = 8'h00;
    ff_ram[7716] = 8'h00;
    ff_ram[7717] = 8'h00;
    ff_ram[7718] = 8'h00;
    ff_ram[7719] = 8'h00;
    ff_ram[7720] = 8'h00;
    ff_ram[7721] = 8'h00;
    ff_ram[7722] = 8'h00;
    ff_ram[7723] = 8'h00;
    ff_ram[7724] = 8'h00;
    ff_ram[7725] = 8'h00;
    ff_ram[7726] = 8'h00;
    ff_ram[7727] = 8'h00;
    ff_ram[7728] = 8'h00;
    ff_ram[7729] = 8'h00;
    ff_ram[7730] = 8'h00;
    ff_ram[7731] = 8'h00;
    ff_ram[7732] = 8'h00;
    ff_ram[7733] = 8'h00;
    ff_ram[7734] = 8'h00;
    ff_ram[7735] = 8'h00;
    ff_ram[7736] = 8'h00;
    ff_ram[7737] = 8'h00;
    ff_ram[7738] = 8'h00;
    ff_ram[7739] = 8'h00;
    ff_ram[7740] = 8'h00;
    ff_ram[7741] = 8'h00;
    ff_ram[7742] = 8'h00;
    ff_ram[7743] = 8'h00;
    ff_ram[7744] = 8'h00;
    ff_ram[7745] = 8'h00;
    ff_ram[7746] = 8'h00;
    ff_ram[7747] = 8'h00;
    ff_ram[7748] = 8'h00;
    ff_ram[7749] = 8'h00;
    ff_ram[7750] = 8'h00;
    ff_ram[7751] = 8'h00;
    ff_ram[7752] = 8'h00;
    ff_ram[7753] = 8'h00;
    ff_ram[7754] = 8'h00;
    ff_ram[7755] = 8'h00;
    ff_ram[7756] = 8'h00;
    ff_ram[7757] = 8'h00;
    ff_ram[7758] = 8'h00;
    ff_ram[7759] = 8'h00;
    ff_ram[7760] = 8'h00;
    ff_ram[7761] = 8'h00;
    ff_ram[7762] = 8'h00;
    ff_ram[7763] = 8'h00;
    ff_ram[7764] = 8'h00;
    ff_ram[7765] = 8'h00;
    ff_ram[7766] = 8'h00;
    ff_ram[7767] = 8'h00;
    ff_ram[7768] = 8'h00;
    ff_ram[7769] = 8'h00;
    ff_ram[7770] = 8'h00;
    ff_ram[7771] = 8'h00;
    ff_ram[7772] = 8'h00;
    ff_ram[7773] = 8'h00;
    ff_ram[7774] = 8'h00;
    ff_ram[7775] = 8'h00;
    ff_ram[7776] = 8'h00;
    ff_ram[7777] = 8'h00;
    ff_ram[7778] = 8'h00;
    ff_ram[7779] = 8'h00;
    ff_ram[7780] = 8'h00;
    ff_ram[7781] = 8'h00;
    ff_ram[7782] = 8'h00;
    ff_ram[7783] = 8'h00;
    ff_ram[7784] = 8'h00;
    ff_ram[7785] = 8'h00;
    ff_ram[7786] = 8'h00;
    ff_ram[7787] = 8'h00;
    ff_ram[7788] = 8'h00;
    ff_ram[7789] = 8'h00;
    ff_ram[7790] = 8'h00;
    ff_ram[7791] = 8'h00;
    ff_ram[7792] = 8'h00;
    ff_ram[7793] = 8'h00;
    ff_ram[7794] = 8'h00;
    ff_ram[7795] = 8'h00;
    ff_ram[7796] = 8'h00;
    ff_ram[7797] = 8'h00;
    ff_ram[7798] = 8'h00;
    ff_ram[7799] = 8'h00;
    ff_ram[7800] = 8'h00;
    ff_ram[7801] = 8'h00;
    ff_ram[7802] = 8'h00;
    ff_ram[7803] = 8'h00;
    ff_ram[7804] = 8'h00;
    ff_ram[7805] = 8'h00;
    ff_ram[7806] = 8'h00;
    ff_ram[7807] = 8'h00;
    ff_ram[7808] = 8'h00;
    ff_ram[7809] = 8'h00;
    ff_ram[7810] = 8'h00;
    ff_ram[7811] = 8'h00;
    ff_ram[7812] = 8'h00;
    ff_ram[7813] = 8'h00;
    ff_ram[7814] = 8'h00;
    ff_ram[7815] = 8'h00;
    ff_ram[7816] = 8'h00;
    ff_ram[7817] = 8'h00;
    ff_ram[7818] = 8'h00;
    ff_ram[7819] = 8'h00;
    ff_ram[7820] = 8'h00;
    ff_ram[7821] = 8'h00;
    ff_ram[7822] = 8'h00;
    ff_ram[7823] = 8'h00;
    ff_ram[7824] = 8'h00;
    ff_ram[7825] = 8'h00;
    ff_ram[7826] = 8'h00;
    ff_ram[7827] = 8'h00;
    ff_ram[7828] = 8'h00;
    ff_ram[7829] = 8'h00;
    ff_ram[7830] = 8'h00;
    ff_ram[7831] = 8'h00;
    ff_ram[7832] = 8'h00;
    ff_ram[7833] = 8'h00;
    ff_ram[7834] = 8'h00;
    ff_ram[7835] = 8'h00;
    ff_ram[7836] = 8'h00;
    ff_ram[7837] = 8'h00;
    ff_ram[7838] = 8'h00;
    ff_ram[7839] = 8'h00;
    ff_ram[7840] = 8'h00;
    ff_ram[7841] = 8'h00;
    ff_ram[7842] = 8'h00;
    ff_ram[7843] = 8'h00;
    ff_ram[7844] = 8'h00;
    ff_ram[7845] = 8'h00;
    ff_ram[7846] = 8'h00;
    ff_ram[7847] = 8'h00;
    ff_ram[7848] = 8'h00;
    ff_ram[7849] = 8'h00;
    ff_ram[7850] = 8'h00;
    ff_ram[7851] = 8'h00;
    ff_ram[7852] = 8'h00;
    ff_ram[7853] = 8'h00;
    ff_ram[7854] = 8'h00;
    ff_ram[7855] = 8'h00;
    ff_ram[7856] = 8'h00;
    ff_ram[7857] = 8'h00;
    ff_ram[7858] = 8'h00;
    ff_ram[7859] = 8'h00;
    ff_ram[7860] = 8'h00;
    ff_ram[7861] = 8'h00;
    ff_ram[7862] = 8'h00;
    ff_ram[7863] = 8'h00;
    ff_ram[7864] = 8'h00;
    ff_ram[7865] = 8'h00;
    ff_ram[7866] = 8'h00;
    ff_ram[7867] = 8'h00;
    ff_ram[7868] = 8'h00;
    ff_ram[7869] = 8'h00;
    ff_ram[7870] = 8'h00;
    ff_ram[7871] = 8'h00;
    ff_ram[7872] = 8'h00;
    ff_ram[7873] = 8'h00;
    ff_ram[7874] = 8'h00;
    ff_ram[7875] = 8'h00;
    ff_ram[7876] = 8'h00;
    ff_ram[7877] = 8'h00;
    ff_ram[7878] = 8'h00;
    ff_ram[7879] = 8'h00;
    ff_ram[7880] = 8'h00;
    ff_ram[7881] = 8'h00;
    ff_ram[7882] = 8'h00;
    ff_ram[7883] = 8'h00;
    ff_ram[7884] = 8'h00;
    ff_ram[7885] = 8'h00;
    ff_ram[7886] = 8'h00;
    ff_ram[7887] = 8'h00;
    ff_ram[7888] = 8'h00;
    ff_ram[7889] = 8'h00;
    ff_ram[7890] = 8'h00;
    ff_ram[7891] = 8'h00;
    ff_ram[7892] = 8'h00;
    ff_ram[7893] = 8'h00;
    ff_ram[7894] = 8'h00;
    ff_ram[7895] = 8'h00;
    ff_ram[7896] = 8'h00;
    ff_ram[7897] = 8'h00;
    ff_ram[7898] = 8'h00;
    ff_ram[7899] = 8'h00;
    ff_ram[7900] = 8'h00;
    ff_ram[7901] = 8'h00;
    ff_ram[7902] = 8'h00;
    ff_ram[7903] = 8'h00;
    ff_ram[7904] = 8'h00;
    ff_ram[7905] = 8'h00;
    ff_ram[7906] = 8'h00;
    ff_ram[7907] = 8'h00;
    ff_ram[7908] = 8'h00;
    ff_ram[7909] = 8'h00;
    ff_ram[7910] = 8'h00;
    ff_ram[7911] = 8'h00;
    ff_ram[7912] = 8'h00;
    ff_ram[7913] = 8'h00;
    ff_ram[7914] = 8'h00;
    ff_ram[7915] = 8'h00;
    ff_ram[7916] = 8'h00;
    ff_ram[7917] = 8'h00;
    ff_ram[7918] = 8'h00;
    ff_ram[7919] = 8'h00;
    ff_ram[7920] = 8'h00;
    ff_ram[7921] = 8'h00;
    ff_ram[7922] = 8'h00;
    ff_ram[7923] = 8'h00;
    ff_ram[7924] = 8'h00;
    ff_ram[7925] = 8'h00;
    ff_ram[7926] = 8'h00;
    ff_ram[7927] = 8'h00;
    ff_ram[7928] = 8'h00;
    ff_ram[7929] = 8'h00;
    ff_ram[7930] = 8'h00;
    ff_ram[7931] = 8'h00;
    ff_ram[7932] = 8'h00;
    ff_ram[7933] = 8'h00;
    ff_ram[7934] = 8'h00;
    ff_ram[7935] = 8'h00;
    ff_ram[7936] = 8'h00;
    ff_ram[7937] = 8'h00;
    ff_ram[7938] = 8'h00;
    ff_ram[7939] = 8'h00;
    ff_ram[7940] = 8'h00;
    ff_ram[7941] = 8'h00;
    ff_ram[7942] = 8'h00;
    ff_ram[7943] = 8'h00;
    ff_ram[7944] = 8'h00;
    ff_ram[7945] = 8'h00;
    ff_ram[7946] = 8'h00;
    ff_ram[7947] = 8'h00;
    ff_ram[7948] = 8'h00;
    ff_ram[7949] = 8'h00;
    ff_ram[7950] = 8'h00;
    ff_ram[7951] = 8'h00;
    ff_ram[7952] = 8'h00;
    ff_ram[7953] = 8'h00;
    ff_ram[7954] = 8'h00;
    ff_ram[7955] = 8'h00;
    ff_ram[7956] = 8'h00;
    ff_ram[7957] = 8'h00;
    ff_ram[7958] = 8'h00;
    ff_ram[7959] = 8'h00;
    ff_ram[7960] = 8'h00;
    ff_ram[7961] = 8'h00;
    ff_ram[7962] = 8'h00;
    ff_ram[7963] = 8'h00;
    ff_ram[7964] = 8'h00;
    ff_ram[7965] = 8'h00;
    ff_ram[7966] = 8'h00;
    ff_ram[7967] = 8'h00;
    ff_ram[7968] = 8'h00;
    ff_ram[7969] = 8'h00;
    ff_ram[7970] = 8'h00;
    ff_ram[7971] = 8'h00;
    ff_ram[7972] = 8'h00;
    ff_ram[7973] = 8'h00;
    ff_ram[7974] = 8'h00;
    ff_ram[7975] = 8'h00;
    ff_ram[7976] = 8'h00;
    ff_ram[7977] = 8'h00;
    ff_ram[7978] = 8'h00;
    ff_ram[7979] = 8'h00;
    ff_ram[7980] = 8'h00;
    ff_ram[7981] = 8'h00;
    ff_ram[7982] = 8'h00;
    ff_ram[7983] = 8'h00;
    ff_ram[7984] = 8'h00;
    ff_ram[7985] = 8'h00;
    ff_ram[7986] = 8'h00;
    ff_ram[7987] = 8'h00;
    ff_ram[7988] = 8'h00;
    ff_ram[7989] = 8'h00;
    ff_ram[7990] = 8'h00;
    ff_ram[7991] = 8'h00;
    ff_ram[7992] = 8'h00;
    ff_ram[7993] = 8'h00;
    ff_ram[7994] = 8'h00;
    ff_ram[7995] = 8'h00;
    ff_ram[7996] = 8'h00;
    ff_ram[7997] = 8'h00;
    ff_ram[7998] = 8'h00;
    ff_ram[7999] = 8'h00;
    ff_ram[8000] = 8'h00;
    ff_ram[8001] = 8'h00;
    ff_ram[8002] = 8'h00;
    ff_ram[8003] = 8'h00;
    ff_ram[8004] = 8'h00;
    ff_ram[8005] = 8'h00;
    ff_ram[8006] = 8'h00;
    ff_ram[8007] = 8'h00;
    ff_ram[8008] = 8'h00;
    ff_ram[8009] = 8'h00;
    ff_ram[8010] = 8'h00;
    ff_ram[8011] = 8'h00;
    ff_ram[8012] = 8'h00;
    ff_ram[8013] = 8'h00;
    ff_ram[8014] = 8'h00;
    ff_ram[8015] = 8'h00;
    ff_ram[8016] = 8'h00;
    ff_ram[8017] = 8'h00;
    ff_ram[8018] = 8'h00;
    ff_ram[8019] = 8'h00;
    ff_ram[8020] = 8'h00;
    ff_ram[8021] = 8'h00;
    ff_ram[8022] = 8'h00;
    ff_ram[8023] = 8'h00;
    ff_ram[8024] = 8'h00;
    ff_ram[8025] = 8'h00;
    ff_ram[8026] = 8'h00;
    ff_ram[8027] = 8'h00;
    ff_ram[8028] = 8'h00;
    ff_ram[8029] = 8'h00;
    ff_ram[8030] = 8'h00;
    ff_ram[8031] = 8'h00;
    ff_ram[8032] = 8'h00;
    ff_ram[8033] = 8'h00;
    ff_ram[8034] = 8'h00;
    ff_ram[8035] = 8'h00;
    ff_ram[8036] = 8'h00;
    ff_ram[8037] = 8'h00;
    ff_ram[8038] = 8'h00;
    ff_ram[8039] = 8'h00;
    ff_ram[8040] = 8'h00;
    ff_ram[8041] = 8'h00;
    ff_ram[8042] = 8'h00;
    ff_ram[8043] = 8'h00;
    ff_ram[8044] = 8'h00;
    ff_ram[8045] = 8'h00;
    ff_ram[8046] = 8'h00;
    ff_ram[8047] = 8'h00;
    ff_ram[8048] = 8'h00;
    ff_ram[8049] = 8'h00;
    ff_ram[8050] = 8'h00;
    ff_ram[8051] = 8'h00;
    ff_ram[8052] = 8'h00;
    ff_ram[8053] = 8'h00;
    ff_ram[8054] = 8'h00;
    ff_ram[8055] = 8'h00;
    ff_ram[8056] = 8'h00;
    ff_ram[8057] = 8'h00;
    ff_ram[8058] = 8'h00;
    ff_ram[8059] = 8'h00;
    ff_ram[8060] = 8'h00;
    ff_ram[8061] = 8'h00;
    ff_ram[8062] = 8'h00;
    ff_ram[8063] = 8'h00;
    ff_ram[8064] = 8'h00;
    ff_ram[8065] = 8'h00;
    ff_ram[8066] = 8'h00;
    ff_ram[8067] = 8'h00;
    ff_ram[8068] = 8'h00;
    ff_ram[8069] = 8'h00;
    ff_ram[8070] = 8'h00;
    ff_ram[8071] = 8'h00;
    ff_ram[8072] = 8'h00;
    ff_ram[8073] = 8'h00;
    ff_ram[8074] = 8'h00;
    ff_ram[8075] = 8'h00;
    ff_ram[8076] = 8'h00;
    ff_ram[8077] = 8'h00;
    ff_ram[8078] = 8'h00;
    ff_ram[8079] = 8'h00;
    ff_ram[8080] = 8'h00;
    ff_ram[8081] = 8'h00;
    ff_ram[8082] = 8'h00;
    ff_ram[8083] = 8'h00;
    ff_ram[8084] = 8'h00;
    ff_ram[8085] = 8'h00;
    ff_ram[8086] = 8'h00;
    ff_ram[8087] = 8'h00;
    ff_ram[8088] = 8'h00;
    ff_ram[8089] = 8'h00;
    ff_ram[8090] = 8'h00;
    ff_ram[8091] = 8'h00;
    ff_ram[8092] = 8'h00;
    ff_ram[8093] = 8'h00;
    ff_ram[8094] = 8'h00;
    ff_ram[8095] = 8'h00;
    ff_ram[8096] = 8'h00;
    ff_ram[8097] = 8'h00;
    ff_ram[8098] = 8'h00;
    ff_ram[8099] = 8'h00;
    ff_ram[8100] = 8'h00;
    ff_ram[8101] = 8'h00;
    ff_ram[8102] = 8'h00;
    ff_ram[8103] = 8'h00;
    ff_ram[8104] = 8'h00;
    ff_ram[8105] = 8'h00;
    ff_ram[8106] = 8'h00;
    ff_ram[8107] = 8'h00;
    ff_ram[8108] = 8'h00;
    ff_ram[8109] = 8'h00;
    ff_ram[8110] = 8'h00;
    ff_ram[8111] = 8'h00;
    ff_ram[8112] = 8'h00;
    ff_ram[8113] = 8'h00;
    ff_ram[8114] = 8'h00;
    ff_ram[8115] = 8'h00;
    ff_ram[8116] = 8'h00;
    ff_ram[8117] = 8'h00;
    ff_ram[8118] = 8'h00;
    ff_ram[8119] = 8'h00;
    ff_ram[8120] = 8'h00;
    ff_ram[8121] = 8'h00;
    ff_ram[8122] = 8'h00;
    ff_ram[8123] = 8'h00;
    ff_ram[8124] = 8'h00;
    ff_ram[8125] = 8'h00;
    ff_ram[8126] = 8'h00;
    ff_ram[8127] = 8'h00;
    ff_ram[8128] = 8'h00;
    ff_ram[8129] = 8'h00;
    ff_ram[8130] = 8'h00;
    ff_ram[8131] = 8'h00;
    ff_ram[8132] = 8'h00;
    ff_ram[8133] = 8'h00;
    ff_ram[8134] = 8'h00;
    ff_ram[8135] = 8'h00;
    ff_ram[8136] = 8'h00;
    ff_ram[8137] = 8'h00;
    ff_ram[8138] = 8'h00;
    ff_ram[8139] = 8'h00;
    ff_ram[8140] = 8'h00;
    ff_ram[8141] = 8'h00;
    ff_ram[8142] = 8'h00;
    ff_ram[8143] = 8'h00;
    ff_ram[8144] = 8'h00;
    ff_ram[8145] = 8'h00;
    ff_ram[8146] = 8'h00;
    ff_ram[8147] = 8'h00;
    ff_ram[8148] = 8'h00;
    ff_ram[8149] = 8'h00;
    ff_ram[8150] = 8'h00;
    ff_ram[8151] = 8'h00;
    ff_ram[8152] = 8'h00;
    ff_ram[8153] = 8'h00;
    ff_ram[8154] = 8'h00;
    ff_ram[8155] = 8'h00;
    ff_ram[8156] = 8'h00;
    ff_ram[8157] = 8'h00;
    ff_ram[8158] = 8'h00;
    ff_ram[8159] = 8'h00;
    ff_ram[8160] = 8'h00;
    ff_ram[8161] = 8'h00;
    ff_ram[8162] = 8'h00;
    ff_ram[8163] = 8'h00;
    ff_ram[8164] = 8'h00;
    ff_ram[8165] = 8'h00;
    ff_ram[8166] = 8'h00;
    ff_ram[8167] = 8'h00;
    ff_ram[8168] = 8'h00;
    ff_ram[8169] = 8'h00;
    ff_ram[8170] = 8'h00;
    ff_ram[8171] = 8'h00;
    ff_ram[8172] = 8'h00;
    ff_ram[8173] = 8'h00;
    ff_ram[8174] = 8'h00;
    ff_ram[8175] = 8'h00;
    ff_ram[8176] = 8'h00;
    ff_ram[8177] = 8'h00;
    ff_ram[8178] = 8'h00;
    ff_ram[8179] = 8'h00;
    ff_ram[8180] = 8'h00;
    ff_ram[8181] = 8'h00;
    ff_ram[8182] = 8'h00;
    ff_ram[8183] = 8'h00;
    ff_ram[8184] = 8'h00;
    ff_ram[8185] = 8'h00;
    ff_ram[8186] = 8'h00;
    ff_ram[8187] = 8'h00;
    ff_ram[8188] = 8'h00;
    ff_ram[8189] = 8'h00;
    ff_ram[8190] = 8'h00;
    ff_ram[8191] = 8'h00;
    ff_ram[8192] = 8'hF4;
    ff_ram[8193] = 8'hF4;
    ff_ram[8194] = 8'hF4;
    ff_ram[8195] = 8'hF4;
    ff_ram[8196] = 8'hF4;
    ff_ram[8197] = 8'hF4;
    ff_ram[8198] = 8'hF4;
    ff_ram[8199] = 8'hF4;
    ff_ram[8200] = 8'hF4;
    ff_ram[8201] = 8'hF4;
    ff_ram[8202] = 8'hF4;
    ff_ram[8203] = 8'hF4;
    ff_ram[8204] = 8'hF4;
    ff_ram[8205] = 8'hF4;
    ff_ram[8206] = 8'hF4;
    ff_ram[8207] = 8'hF4;
    ff_ram[8208] = 8'hF4;
    ff_ram[8209] = 8'hF4;
    ff_ram[8210] = 8'hF4;
    ff_ram[8211] = 8'hF4;
    ff_ram[8212] = 8'hF4;
    ff_ram[8213] = 8'hF4;
    ff_ram[8214] = 8'hF4;
    ff_ram[8215] = 8'hF4;
    ff_ram[8216] = 8'hF4;
    ff_ram[8217] = 8'hF4;
    ff_ram[8218] = 8'hF4;
    ff_ram[8219] = 8'hF4;
    ff_ram[8220] = 8'hF4;
    ff_ram[8221] = 8'hF4;
    ff_ram[8222] = 8'hF4;
    ff_ram[8223] = 8'hF4;
    ff_ram[8224] = 8'h00;
    ff_ram[8225] = 8'h00;
    ff_ram[8226] = 8'h00;
    ff_ram[8227] = 8'h00;
    ff_ram[8228] = 8'h11;
    ff_ram[8229] = 8'h06;
    ff_ram[8230] = 8'h33;
    ff_ram[8231] = 8'h07;
    ff_ram[8232] = 8'h17;
    ff_ram[8233] = 8'h01;
    ff_ram[8234] = 8'h27;
    ff_ram[8235] = 8'h03;
    ff_ram[8236] = 8'h51;
    ff_ram[8237] = 8'h01;
    ff_ram[8238] = 8'h27;
    ff_ram[8239] = 8'h06;
    ff_ram[8240] = 8'h71;
    ff_ram[8241] = 8'h01;
    ff_ram[8242] = 8'h73;
    ff_ram[8243] = 8'h03;
    ff_ram[8244] = 8'h61;
    ff_ram[8245] = 8'h06;
    ff_ram[8246] = 8'h64;
    ff_ram[8247] = 8'h06;
    ff_ram[8248] = 8'h11;
    ff_ram[8249] = 8'h04;
    ff_ram[8250] = 8'h65;
    ff_ram[8251] = 8'h02;
    ff_ram[8252] = 8'h55;
    ff_ram[8253] = 8'h05;
    ff_ram[8254] = 8'h77;
    ff_ram[8255] = 8'h07;
    ff_ram[8256] = 8'h00;
    ff_ram[8257] = 8'h00;
    ff_ram[8258] = 8'h00;
    ff_ram[8259] = 8'h00;
    ff_ram[8260] = 8'h00;
    ff_ram[8261] = 8'h00;
    ff_ram[8262] = 8'h00;
    ff_ram[8263] = 8'h00;
    ff_ram[8264] = 8'h00;
    ff_ram[8265] = 8'h00;
    ff_ram[8266] = 8'h00;
    ff_ram[8267] = 8'h00;
    ff_ram[8268] = 8'h00;
    ff_ram[8269] = 8'h00;
    ff_ram[8270] = 8'h00;
    ff_ram[8271] = 8'h00;
    ff_ram[8272] = 8'h00;
    ff_ram[8273] = 8'h00;
    ff_ram[8274] = 8'h00;
    ff_ram[8275] = 8'h00;
    ff_ram[8276] = 8'h00;
    ff_ram[8277] = 8'h00;
    ff_ram[8278] = 8'h00;
    ff_ram[8279] = 8'h00;
    ff_ram[8280] = 8'h00;
    ff_ram[8281] = 8'h00;
    ff_ram[8282] = 8'h00;
    ff_ram[8283] = 8'h00;
    ff_ram[8284] = 8'h00;
    ff_ram[8285] = 8'h00;
    ff_ram[8286] = 8'h00;
    ff_ram[8287] = 8'h00;
    ff_ram[8288] = 8'h00;
    ff_ram[8289] = 8'h00;
    ff_ram[8290] = 8'h00;
    ff_ram[8291] = 8'h00;
    ff_ram[8292] = 8'h00;
    ff_ram[8293] = 8'h00;
    ff_ram[8294] = 8'h00;
    ff_ram[8295] = 8'h00;
    ff_ram[8296] = 8'h00;
    ff_ram[8297] = 8'h00;
    ff_ram[8298] = 8'h00;
    ff_ram[8299] = 8'h00;
    ff_ram[8300] = 8'h00;
    ff_ram[8301] = 8'h00;
    ff_ram[8302] = 8'h00;
    ff_ram[8303] = 8'h00;
    ff_ram[8304] = 8'h00;
    ff_ram[8305] = 8'h00;
    ff_ram[8306] = 8'h00;
    ff_ram[8307] = 8'h00;
    ff_ram[8308] = 8'h00;
    ff_ram[8309] = 8'h00;
    ff_ram[8310] = 8'h00;
    ff_ram[8311] = 8'h00;
    ff_ram[8312] = 8'h00;
    ff_ram[8313] = 8'h00;
    ff_ram[8314] = 8'h00;
    ff_ram[8315] = 8'h00;
    ff_ram[8316] = 8'h00;
    ff_ram[8317] = 8'h00;
    ff_ram[8318] = 8'h00;
    ff_ram[8319] = 8'h00;
    ff_ram[8320] = 8'h00;
    ff_ram[8321] = 8'h00;
    ff_ram[8322] = 8'h00;
    ff_ram[8323] = 8'h00;
    ff_ram[8324] = 8'h00;
    ff_ram[8325] = 8'h00;
    ff_ram[8326] = 8'h00;
    ff_ram[8327] = 8'h00;
    ff_ram[8328] = 8'h00;
    ff_ram[8329] = 8'h00;
    ff_ram[8330] = 8'h00;
    ff_ram[8331] = 8'h00;
    ff_ram[8332] = 8'h00;
    ff_ram[8333] = 8'h00;
    ff_ram[8334] = 8'h00;
    ff_ram[8335] = 8'h00;
    ff_ram[8336] = 8'h00;
    ff_ram[8337] = 8'h00;
    ff_ram[8338] = 8'h00;
    ff_ram[8339] = 8'h00;
    ff_ram[8340] = 8'h00;
    ff_ram[8341] = 8'h00;
    ff_ram[8342] = 8'h00;
    ff_ram[8343] = 8'h00;
    ff_ram[8344] = 8'h00;
    ff_ram[8345] = 8'h00;
    ff_ram[8346] = 8'h00;
    ff_ram[8347] = 8'h00;
    ff_ram[8348] = 8'h00;
    ff_ram[8349] = 8'h00;
    ff_ram[8350] = 8'h00;
    ff_ram[8351] = 8'h00;
    ff_ram[8352] = 8'h00;
    ff_ram[8353] = 8'h00;
    ff_ram[8354] = 8'h00;
    ff_ram[8355] = 8'h00;
    ff_ram[8356] = 8'h00;
    ff_ram[8357] = 8'h00;
    ff_ram[8358] = 8'h00;
    ff_ram[8359] = 8'h00;
    ff_ram[8360] = 8'h00;
    ff_ram[8361] = 8'h00;
    ff_ram[8362] = 8'h00;
    ff_ram[8363] = 8'h00;
    ff_ram[8364] = 8'h00;
    ff_ram[8365] = 8'h00;
    ff_ram[8366] = 8'h00;
    ff_ram[8367] = 8'h00;
    ff_ram[8368] = 8'h00;
    ff_ram[8369] = 8'h00;
    ff_ram[8370] = 8'h00;
    ff_ram[8371] = 8'h00;
    ff_ram[8372] = 8'h00;
    ff_ram[8373] = 8'h00;
    ff_ram[8374] = 8'h00;
    ff_ram[8375] = 8'h00;
    ff_ram[8376] = 8'h00;
    ff_ram[8377] = 8'h00;
    ff_ram[8378] = 8'h00;
    ff_ram[8379] = 8'h00;
    ff_ram[8380] = 8'h00;
    ff_ram[8381] = 8'h00;
    ff_ram[8382] = 8'h00;
    ff_ram[8383] = 8'h00;
    ff_ram[8384] = 8'h00;
    ff_ram[8385] = 8'h00;
    ff_ram[8386] = 8'h00;
    ff_ram[8387] = 8'h00;
    ff_ram[8388] = 8'h00;
    ff_ram[8389] = 8'h00;
    ff_ram[8390] = 8'h00;
    ff_ram[8391] = 8'h00;
    ff_ram[8392] = 8'h00;
    ff_ram[8393] = 8'h00;
    ff_ram[8394] = 8'h00;
    ff_ram[8395] = 8'h00;
    ff_ram[8396] = 8'h00;
    ff_ram[8397] = 8'h00;
    ff_ram[8398] = 8'h00;
    ff_ram[8399] = 8'h00;
    ff_ram[8400] = 8'h00;
    ff_ram[8401] = 8'h00;
    ff_ram[8402] = 8'h00;
    ff_ram[8403] = 8'h00;
    ff_ram[8404] = 8'h00;
    ff_ram[8405] = 8'h00;
    ff_ram[8406] = 8'h00;
    ff_ram[8407] = 8'h00;
    ff_ram[8408] = 8'h00;
    ff_ram[8409] = 8'h00;
    ff_ram[8410] = 8'h00;
    ff_ram[8411] = 8'h00;
    ff_ram[8412] = 8'h00;
    ff_ram[8413] = 8'h00;
    ff_ram[8414] = 8'h00;
    ff_ram[8415] = 8'h00;
    ff_ram[8416] = 8'h00;
    ff_ram[8417] = 8'h00;
    ff_ram[8418] = 8'h00;
    ff_ram[8419] = 8'h00;
    ff_ram[8420] = 8'h00;
    ff_ram[8421] = 8'h00;
    ff_ram[8422] = 8'h00;
    ff_ram[8423] = 8'h00;
    ff_ram[8424] = 8'h00;
    ff_ram[8425] = 8'h00;
    ff_ram[8426] = 8'h00;
    ff_ram[8427] = 8'h00;
    ff_ram[8428] = 8'h00;
    ff_ram[8429] = 8'h00;
    ff_ram[8430] = 8'h00;
    ff_ram[8431] = 8'h00;
    ff_ram[8432] = 8'h00;
    ff_ram[8433] = 8'h00;
    ff_ram[8434] = 8'h00;
    ff_ram[8435] = 8'h00;
    ff_ram[8436] = 8'h00;
    ff_ram[8437] = 8'h00;
    ff_ram[8438] = 8'h00;
    ff_ram[8439] = 8'h00;
    ff_ram[8440] = 8'h00;
    ff_ram[8441] = 8'h00;
    ff_ram[8442] = 8'h00;
    ff_ram[8443] = 8'h00;
    ff_ram[8444] = 8'h00;
    ff_ram[8445] = 8'h00;
    ff_ram[8446] = 8'h00;
    ff_ram[8447] = 8'h00;
    ff_ram[8448] = 8'h00;
    ff_ram[8449] = 8'h00;
    ff_ram[8450] = 8'h00;
    ff_ram[8451] = 8'h00;
    ff_ram[8452] = 8'h00;
    ff_ram[8453] = 8'h00;
    ff_ram[8454] = 8'h00;
    ff_ram[8455] = 8'h00;
    ff_ram[8456] = 8'h00;
    ff_ram[8457] = 8'h00;
    ff_ram[8458] = 8'h00;
    ff_ram[8459] = 8'h00;
    ff_ram[8460] = 8'h00;
    ff_ram[8461] = 8'h00;
    ff_ram[8462] = 8'h00;
    ff_ram[8463] = 8'h00;
    ff_ram[8464] = 8'h00;
    ff_ram[8465] = 8'h00;
    ff_ram[8466] = 8'h00;
    ff_ram[8467] = 8'h00;
    ff_ram[8468] = 8'h00;
    ff_ram[8469] = 8'h00;
    ff_ram[8470] = 8'h00;
    ff_ram[8471] = 8'h00;
    ff_ram[8472] = 8'h00;
    ff_ram[8473] = 8'h00;
    ff_ram[8474] = 8'h00;
    ff_ram[8475] = 8'h00;
    ff_ram[8476] = 8'h00;
    ff_ram[8477] = 8'h00;
    ff_ram[8478] = 8'h00;
    ff_ram[8479] = 8'h00;
    ff_ram[8480] = 8'h00;
    ff_ram[8481] = 8'h00;
    ff_ram[8482] = 8'h00;
    ff_ram[8483] = 8'h00;
    ff_ram[8484] = 8'h00;
    ff_ram[8485] = 8'h00;
    ff_ram[8486] = 8'h00;
    ff_ram[8487] = 8'h00;
    ff_ram[8488] = 8'h00;
    ff_ram[8489] = 8'h00;
    ff_ram[8490] = 8'h00;
    ff_ram[8491] = 8'h00;
    ff_ram[8492] = 8'h00;
    ff_ram[8493] = 8'h00;
    ff_ram[8494] = 8'h00;
    ff_ram[8495] = 8'h00;
    ff_ram[8496] = 8'h00;
    ff_ram[8497] = 8'h00;
    ff_ram[8498] = 8'h00;
    ff_ram[8499] = 8'h00;
    ff_ram[8500] = 8'h00;
    ff_ram[8501] = 8'h00;
    ff_ram[8502] = 8'h00;
    ff_ram[8503] = 8'h00;
    ff_ram[8504] = 8'h00;
    ff_ram[8505] = 8'h00;
    ff_ram[8506] = 8'h00;
    ff_ram[8507] = 8'h00;
    ff_ram[8508] = 8'h00;
    ff_ram[8509] = 8'h00;
    ff_ram[8510] = 8'h00;
    ff_ram[8511] = 8'h00;
    ff_ram[8512] = 8'h00;
    ff_ram[8513] = 8'h00;
    ff_ram[8514] = 8'h00;
    ff_ram[8515] = 8'h00;
    ff_ram[8516] = 8'h00;
    ff_ram[8517] = 8'h00;
    ff_ram[8518] = 8'h00;
    ff_ram[8519] = 8'h00;
    ff_ram[8520] = 8'h00;
    ff_ram[8521] = 8'h00;
    ff_ram[8522] = 8'h00;
    ff_ram[8523] = 8'h00;
    ff_ram[8524] = 8'h00;
    ff_ram[8525] = 8'h00;
    ff_ram[8526] = 8'h00;
    ff_ram[8527] = 8'h00;
    ff_ram[8528] = 8'h00;
    ff_ram[8529] = 8'h00;
    ff_ram[8530] = 8'h00;
    ff_ram[8531] = 8'h00;
    ff_ram[8532] = 8'h00;
    ff_ram[8533] = 8'h00;
    ff_ram[8534] = 8'h00;
    ff_ram[8535] = 8'h00;
    ff_ram[8536] = 8'h00;
    ff_ram[8537] = 8'h00;
    ff_ram[8538] = 8'h00;
    ff_ram[8539] = 8'h00;
    ff_ram[8540] = 8'h00;
    ff_ram[8541] = 8'h00;
    ff_ram[8542] = 8'h00;
    ff_ram[8543] = 8'h00;
    ff_ram[8544] = 8'h00;
    ff_ram[8545] = 8'h00;
    ff_ram[8546] = 8'h00;
    ff_ram[8547] = 8'h00;
    ff_ram[8548] = 8'h00;
    ff_ram[8549] = 8'h00;
    ff_ram[8550] = 8'h00;
    ff_ram[8551] = 8'h00;
    ff_ram[8552] = 8'h00;
    ff_ram[8553] = 8'h00;
    ff_ram[8554] = 8'h00;
    ff_ram[8555] = 8'h00;
    ff_ram[8556] = 8'h00;
    ff_ram[8557] = 8'h00;
    ff_ram[8558] = 8'h00;
    ff_ram[8559] = 8'h00;
    ff_ram[8560] = 8'h00;
    ff_ram[8561] = 8'h00;
    ff_ram[8562] = 8'h00;
    ff_ram[8563] = 8'h00;
    ff_ram[8564] = 8'h00;
    ff_ram[8565] = 8'h00;
    ff_ram[8566] = 8'h00;
    ff_ram[8567] = 8'h00;
    ff_ram[8568] = 8'h00;
    ff_ram[8569] = 8'h00;
    ff_ram[8570] = 8'h00;
    ff_ram[8571] = 8'h00;
    ff_ram[8572] = 8'h00;
    ff_ram[8573] = 8'h00;
    ff_ram[8574] = 8'h00;
    ff_ram[8575] = 8'h00;
    ff_ram[8576] = 8'h00;
    ff_ram[8577] = 8'h00;
    ff_ram[8578] = 8'h00;
    ff_ram[8579] = 8'h00;
    ff_ram[8580] = 8'h00;
    ff_ram[8581] = 8'h00;
    ff_ram[8582] = 8'h00;
    ff_ram[8583] = 8'h00;
    ff_ram[8584] = 8'h00;
    ff_ram[8585] = 8'h00;
    ff_ram[8586] = 8'h00;
    ff_ram[8587] = 8'h00;
    ff_ram[8588] = 8'h00;
    ff_ram[8589] = 8'h00;
    ff_ram[8590] = 8'h00;
    ff_ram[8591] = 8'h00;
    ff_ram[8592] = 8'h00;
    ff_ram[8593] = 8'h00;
    ff_ram[8594] = 8'h00;
    ff_ram[8595] = 8'h00;
    ff_ram[8596] = 8'h00;
    ff_ram[8597] = 8'h00;
    ff_ram[8598] = 8'h00;
    ff_ram[8599] = 8'h00;
    ff_ram[8600] = 8'h00;
    ff_ram[8601] = 8'h00;
    ff_ram[8602] = 8'h00;
    ff_ram[8603] = 8'h00;
    ff_ram[8604] = 8'h00;
    ff_ram[8605] = 8'h00;
    ff_ram[8606] = 8'h00;
    ff_ram[8607] = 8'h00;
    ff_ram[8608] = 8'h00;
    ff_ram[8609] = 8'h00;
    ff_ram[8610] = 8'h00;
    ff_ram[8611] = 8'h00;
    ff_ram[8612] = 8'h00;
    ff_ram[8613] = 8'h00;
    ff_ram[8614] = 8'h00;
    ff_ram[8615] = 8'h00;
    ff_ram[8616] = 8'h00;
    ff_ram[8617] = 8'h00;
    ff_ram[8618] = 8'h00;
    ff_ram[8619] = 8'h00;
    ff_ram[8620] = 8'h00;
    ff_ram[8621] = 8'h00;
    ff_ram[8622] = 8'h00;
    ff_ram[8623] = 8'h00;
    ff_ram[8624] = 8'h00;
    ff_ram[8625] = 8'h00;
    ff_ram[8626] = 8'h00;
    ff_ram[8627] = 8'h00;
    ff_ram[8628] = 8'h00;
    ff_ram[8629] = 8'h00;
    ff_ram[8630] = 8'h00;
    ff_ram[8631] = 8'h00;
    ff_ram[8632] = 8'h00;
    ff_ram[8633] = 8'h00;
    ff_ram[8634] = 8'h00;
    ff_ram[8635] = 8'h00;
    ff_ram[8636] = 8'h00;
    ff_ram[8637] = 8'h00;
    ff_ram[8638] = 8'h00;
    ff_ram[8639] = 8'h00;
    ff_ram[8640] = 8'h00;
    ff_ram[8641] = 8'h00;
    ff_ram[8642] = 8'h00;
    ff_ram[8643] = 8'h00;
    ff_ram[8644] = 8'h00;
    ff_ram[8645] = 8'h00;
    ff_ram[8646] = 8'h00;
    ff_ram[8647] = 8'h00;
    ff_ram[8648] = 8'h00;
    ff_ram[8649] = 8'h00;
    ff_ram[8650] = 8'h00;
    ff_ram[8651] = 8'h00;
    ff_ram[8652] = 8'h00;
    ff_ram[8653] = 8'h00;
    ff_ram[8654] = 8'h00;
    ff_ram[8655] = 8'h00;
    ff_ram[8656] = 8'h00;
    ff_ram[8657] = 8'h00;
    ff_ram[8658] = 8'h00;
    ff_ram[8659] = 8'h00;
    ff_ram[8660] = 8'h00;
    ff_ram[8661] = 8'h00;
    ff_ram[8662] = 8'h00;
    ff_ram[8663] = 8'h00;
    ff_ram[8664] = 8'h00;
    ff_ram[8665] = 8'h00;
    ff_ram[8666] = 8'h00;
    ff_ram[8667] = 8'h00;
    ff_ram[8668] = 8'h00;
    ff_ram[8669] = 8'h00;
    ff_ram[8670] = 8'h00;
    ff_ram[8671] = 8'h00;
    ff_ram[8672] = 8'h00;
    ff_ram[8673] = 8'h00;
    ff_ram[8674] = 8'h00;
    ff_ram[8675] = 8'h00;
    ff_ram[8676] = 8'h00;
    ff_ram[8677] = 8'h00;
    ff_ram[8678] = 8'h00;
    ff_ram[8679] = 8'h00;
    ff_ram[8680] = 8'h00;
    ff_ram[8681] = 8'h00;
    ff_ram[8682] = 8'h00;
    ff_ram[8683] = 8'h00;
    ff_ram[8684] = 8'h00;
    ff_ram[8685] = 8'h00;
    ff_ram[8686] = 8'h00;
    ff_ram[8687] = 8'h00;
    ff_ram[8688] = 8'h00;
    ff_ram[8689] = 8'h00;
    ff_ram[8690] = 8'h00;
    ff_ram[8691] = 8'h00;
    ff_ram[8692] = 8'h00;
    ff_ram[8693] = 8'h00;
    ff_ram[8694] = 8'h00;
    ff_ram[8695] = 8'h00;
    ff_ram[8696] = 8'h00;
    ff_ram[8697] = 8'h00;
    ff_ram[8698] = 8'h00;
    ff_ram[8699] = 8'h00;
    ff_ram[8700] = 8'h00;
    ff_ram[8701] = 8'h00;
    ff_ram[8702] = 8'h00;
    ff_ram[8703] = 8'h00;
    ff_ram[8704] = 8'h00;
    ff_ram[8705] = 8'h00;
    ff_ram[8706] = 8'h00;
    ff_ram[8707] = 8'h00;
    ff_ram[8708] = 8'h00;
    ff_ram[8709] = 8'h00;
    ff_ram[8710] = 8'h00;
    ff_ram[8711] = 8'h00;
    ff_ram[8712] = 8'h00;
    ff_ram[8713] = 8'h00;
    ff_ram[8714] = 8'h00;
    ff_ram[8715] = 8'h00;
    ff_ram[8716] = 8'h00;
    ff_ram[8717] = 8'h00;
    ff_ram[8718] = 8'h00;
    ff_ram[8719] = 8'h00;
    ff_ram[8720] = 8'h00;
    ff_ram[8721] = 8'h00;
    ff_ram[8722] = 8'h00;
    ff_ram[8723] = 8'h00;
    ff_ram[8724] = 8'h00;
    ff_ram[8725] = 8'h00;
    ff_ram[8726] = 8'h00;
    ff_ram[8727] = 8'h00;
    ff_ram[8728] = 8'h00;
    ff_ram[8729] = 8'h00;
    ff_ram[8730] = 8'h00;
    ff_ram[8731] = 8'h00;
    ff_ram[8732] = 8'h00;
    ff_ram[8733] = 8'h00;
    ff_ram[8734] = 8'h00;
    ff_ram[8735] = 8'h00;
    ff_ram[8736] = 8'h00;
    ff_ram[8737] = 8'h00;
    ff_ram[8738] = 8'h00;
    ff_ram[8739] = 8'h00;
    ff_ram[8740] = 8'h00;
    ff_ram[8741] = 8'h00;
    ff_ram[8742] = 8'h00;
    ff_ram[8743] = 8'h00;
    ff_ram[8744] = 8'h00;
    ff_ram[8745] = 8'h00;
    ff_ram[8746] = 8'h00;
    ff_ram[8747] = 8'h00;
    ff_ram[8748] = 8'h00;
    ff_ram[8749] = 8'h00;
    ff_ram[8750] = 8'h00;
    ff_ram[8751] = 8'h00;
    ff_ram[8752] = 8'h00;
    ff_ram[8753] = 8'h00;
    ff_ram[8754] = 8'h00;
    ff_ram[8755] = 8'h00;
    ff_ram[8756] = 8'h00;
    ff_ram[8757] = 8'h00;
    ff_ram[8758] = 8'h00;
    ff_ram[8759] = 8'h00;
    ff_ram[8760] = 8'h00;
    ff_ram[8761] = 8'h00;
    ff_ram[8762] = 8'h00;
    ff_ram[8763] = 8'h00;
    ff_ram[8764] = 8'h00;
    ff_ram[8765] = 8'h00;
    ff_ram[8766] = 8'h00;
    ff_ram[8767] = 8'h00;
    ff_ram[8768] = 8'h00;
    ff_ram[8769] = 8'h00;
    ff_ram[8770] = 8'h00;
    ff_ram[8771] = 8'h00;
    ff_ram[8772] = 8'h00;
    ff_ram[8773] = 8'h00;
    ff_ram[8774] = 8'h00;
    ff_ram[8775] = 8'h00;
    ff_ram[8776] = 8'h00;
    ff_ram[8777] = 8'h00;
    ff_ram[8778] = 8'h00;
    ff_ram[8779] = 8'h00;
    ff_ram[8780] = 8'h00;
    ff_ram[8781] = 8'h00;
    ff_ram[8782] = 8'h00;
    ff_ram[8783] = 8'h00;
    ff_ram[8784] = 8'h00;
    ff_ram[8785] = 8'h00;
    ff_ram[8786] = 8'h00;
    ff_ram[8787] = 8'h00;
    ff_ram[8788] = 8'h00;
    ff_ram[8789] = 8'h00;
    ff_ram[8790] = 8'h00;
    ff_ram[8791] = 8'h00;
    ff_ram[8792] = 8'h00;
    ff_ram[8793] = 8'h00;
    ff_ram[8794] = 8'h00;
    ff_ram[8795] = 8'h00;
    ff_ram[8796] = 8'h00;
    ff_ram[8797] = 8'h00;
    ff_ram[8798] = 8'h00;
    ff_ram[8799] = 8'h00;
    ff_ram[8800] = 8'h00;
    ff_ram[8801] = 8'h00;
    ff_ram[8802] = 8'h00;
    ff_ram[8803] = 8'h00;
    ff_ram[8804] = 8'h00;
    ff_ram[8805] = 8'h00;
    ff_ram[8806] = 8'h00;
    ff_ram[8807] = 8'h00;
    ff_ram[8808] = 8'h00;
    ff_ram[8809] = 8'h00;
    ff_ram[8810] = 8'h00;
    ff_ram[8811] = 8'h00;
    ff_ram[8812] = 8'h00;
    ff_ram[8813] = 8'h00;
    ff_ram[8814] = 8'h00;
    ff_ram[8815] = 8'h00;
    ff_ram[8816] = 8'h00;
    ff_ram[8817] = 8'h00;
    ff_ram[8818] = 8'h00;
    ff_ram[8819] = 8'h00;
    ff_ram[8820] = 8'h00;
    ff_ram[8821] = 8'h00;
    ff_ram[8822] = 8'h00;
    ff_ram[8823] = 8'h00;
    ff_ram[8824] = 8'h00;
    ff_ram[8825] = 8'h00;
    ff_ram[8826] = 8'h00;
    ff_ram[8827] = 8'h00;
    ff_ram[8828] = 8'h00;
    ff_ram[8829] = 8'h00;
    ff_ram[8830] = 8'h00;
    ff_ram[8831] = 8'h00;
    ff_ram[8832] = 8'h00;
    ff_ram[8833] = 8'h00;
    ff_ram[8834] = 8'h00;
    ff_ram[8835] = 8'h00;
    ff_ram[8836] = 8'h00;
    ff_ram[8837] = 8'h00;
    ff_ram[8838] = 8'h00;
    ff_ram[8839] = 8'h00;
    ff_ram[8840] = 8'h00;
    ff_ram[8841] = 8'h00;
    ff_ram[8842] = 8'h00;
    ff_ram[8843] = 8'h00;
    ff_ram[8844] = 8'h00;
    ff_ram[8845] = 8'h00;
    ff_ram[8846] = 8'h00;
    ff_ram[8847] = 8'h00;
    ff_ram[8848] = 8'h00;
    ff_ram[8849] = 8'h00;
    ff_ram[8850] = 8'h00;
    ff_ram[8851] = 8'h00;
    ff_ram[8852] = 8'h00;
    ff_ram[8853] = 8'h00;
    ff_ram[8854] = 8'h00;
    ff_ram[8855] = 8'h00;
    ff_ram[8856] = 8'h00;
    ff_ram[8857] = 8'h00;
    ff_ram[8858] = 8'h00;
    ff_ram[8859] = 8'h00;
    ff_ram[8860] = 8'h00;
    ff_ram[8861] = 8'h00;
    ff_ram[8862] = 8'h00;
    ff_ram[8863] = 8'h00;
    ff_ram[8864] = 8'h00;
    ff_ram[8865] = 8'h00;
    ff_ram[8866] = 8'h00;
    ff_ram[8867] = 8'h00;
    ff_ram[8868] = 8'h00;
    ff_ram[8869] = 8'h00;
    ff_ram[8870] = 8'h00;
    ff_ram[8871] = 8'h00;
    ff_ram[8872] = 8'h00;
    ff_ram[8873] = 8'h00;
    ff_ram[8874] = 8'h00;
    ff_ram[8875] = 8'h00;
    ff_ram[8876] = 8'h00;
    ff_ram[8877] = 8'h00;
    ff_ram[8878] = 8'h00;
    ff_ram[8879] = 8'h00;
    ff_ram[8880] = 8'h00;
    ff_ram[8881] = 8'h00;
    ff_ram[8882] = 8'h00;
    ff_ram[8883] = 8'h00;
    ff_ram[8884] = 8'h00;
    ff_ram[8885] = 8'h00;
    ff_ram[8886] = 8'h00;
    ff_ram[8887] = 8'h00;
    ff_ram[8888] = 8'h00;
    ff_ram[8889] = 8'h00;
    ff_ram[8890] = 8'h00;
    ff_ram[8891] = 8'h00;
    ff_ram[8892] = 8'h00;
    ff_ram[8893] = 8'h00;
    ff_ram[8894] = 8'h00;
    ff_ram[8895] = 8'h00;
    ff_ram[8896] = 8'h00;
    ff_ram[8897] = 8'h00;
    ff_ram[8898] = 8'h00;
    ff_ram[8899] = 8'h00;
    ff_ram[8900] = 8'h00;
    ff_ram[8901] = 8'h00;
    ff_ram[8902] = 8'h00;
    ff_ram[8903] = 8'h00;
    ff_ram[8904] = 8'h00;
    ff_ram[8905] = 8'h00;
    ff_ram[8906] = 8'h00;
    ff_ram[8907] = 8'h00;
    ff_ram[8908] = 8'h00;
    ff_ram[8909] = 8'h00;
    ff_ram[8910] = 8'h00;
    ff_ram[8911] = 8'h00;
    ff_ram[8912] = 8'h00;
    ff_ram[8913] = 8'h00;
    ff_ram[8914] = 8'h00;
    ff_ram[8915] = 8'h00;
    ff_ram[8916] = 8'h00;
    ff_ram[8917] = 8'h00;
    ff_ram[8918] = 8'h00;
    ff_ram[8919] = 8'h00;
    ff_ram[8920] = 8'h00;
    ff_ram[8921] = 8'h00;
    ff_ram[8922] = 8'h00;
    ff_ram[8923] = 8'h00;
    ff_ram[8924] = 8'h00;
    ff_ram[8925] = 8'h00;
    ff_ram[8926] = 8'h00;
    ff_ram[8927] = 8'h00;
    ff_ram[8928] = 8'h00;
    ff_ram[8929] = 8'h00;
    ff_ram[8930] = 8'h00;
    ff_ram[8931] = 8'h00;
    ff_ram[8932] = 8'h00;
    ff_ram[8933] = 8'h00;
    ff_ram[8934] = 8'h00;
    ff_ram[8935] = 8'h00;
    ff_ram[8936] = 8'h00;
    ff_ram[8937] = 8'h00;
    ff_ram[8938] = 8'h00;
    ff_ram[8939] = 8'h00;
    ff_ram[8940] = 8'h00;
    ff_ram[8941] = 8'h00;
    ff_ram[8942] = 8'h00;
    ff_ram[8943] = 8'h00;
    ff_ram[8944] = 8'h00;
    ff_ram[8945] = 8'h00;
    ff_ram[8946] = 8'h00;
    ff_ram[8947] = 8'h00;
    ff_ram[8948] = 8'h00;
    ff_ram[8949] = 8'h00;
    ff_ram[8950] = 8'h00;
    ff_ram[8951] = 8'h00;
    ff_ram[8952] = 8'h00;
    ff_ram[8953] = 8'h00;
    ff_ram[8954] = 8'h00;
    ff_ram[8955] = 8'h00;
    ff_ram[8956] = 8'h00;
    ff_ram[8957] = 8'h00;
    ff_ram[8958] = 8'h00;
    ff_ram[8959] = 8'h00;
    ff_ram[8960] = 8'h00;
    ff_ram[8961] = 8'h00;
    ff_ram[8962] = 8'h00;
    ff_ram[8963] = 8'h00;
    ff_ram[8964] = 8'h00;
    ff_ram[8965] = 8'h00;
    ff_ram[8966] = 8'h00;
    ff_ram[8967] = 8'h00;
    ff_ram[8968] = 8'h00;
    ff_ram[8969] = 8'h00;
    ff_ram[8970] = 8'h00;
    ff_ram[8971] = 8'h00;
    ff_ram[8972] = 8'h00;
    ff_ram[8973] = 8'h00;
    ff_ram[8974] = 8'h00;
    ff_ram[8975] = 8'h00;
    ff_ram[8976] = 8'h00;
    ff_ram[8977] = 8'h00;
    ff_ram[8978] = 8'h00;
    ff_ram[8979] = 8'h00;
    ff_ram[8980] = 8'h00;
    ff_ram[8981] = 8'h00;
    ff_ram[8982] = 8'h00;
    ff_ram[8983] = 8'h00;
    ff_ram[8984] = 8'h00;
    ff_ram[8985] = 8'h00;
    ff_ram[8986] = 8'h00;
    ff_ram[8987] = 8'h00;
    ff_ram[8988] = 8'h00;
    ff_ram[8989] = 8'h00;
    ff_ram[8990] = 8'h00;
    ff_ram[8991] = 8'h00;
    ff_ram[8992] = 8'h00;
    ff_ram[8993] = 8'h00;
    ff_ram[8994] = 8'h00;
    ff_ram[8995] = 8'h00;
    ff_ram[8996] = 8'h00;
    ff_ram[8997] = 8'h00;
    ff_ram[8998] = 8'h00;
    ff_ram[8999] = 8'h00;
    ff_ram[9000] = 8'h00;
    ff_ram[9001] = 8'h00;
    ff_ram[9002] = 8'h00;
    ff_ram[9003] = 8'h00;
    ff_ram[9004] = 8'h00;
    ff_ram[9005] = 8'h00;
    ff_ram[9006] = 8'h00;
    ff_ram[9007] = 8'h00;
    ff_ram[9008] = 8'h00;
    ff_ram[9009] = 8'h00;
    ff_ram[9010] = 8'h00;
    ff_ram[9011] = 8'h00;
    ff_ram[9012] = 8'h00;
    ff_ram[9013] = 8'h00;
    ff_ram[9014] = 8'h00;
    ff_ram[9015] = 8'h00;
    ff_ram[9016] = 8'h00;
    ff_ram[9017] = 8'h00;
    ff_ram[9018] = 8'h00;
    ff_ram[9019] = 8'h00;
    ff_ram[9020] = 8'h00;
    ff_ram[9021] = 8'h00;
    ff_ram[9022] = 8'h00;
    ff_ram[9023] = 8'h00;
    ff_ram[9024] = 8'h00;
    ff_ram[9025] = 8'h00;
    ff_ram[9026] = 8'h00;
    ff_ram[9027] = 8'h00;
    ff_ram[9028] = 8'h00;
    ff_ram[9029] = 8'h00;
    ff_ram[9030] = 8'h00;
    ff_ram[9031] = 8'h00;
    ff_ram[9032] = 8'h00;
    ff_ram[9033] = 8'h00;
    ff_ram[9034] = 8'h00;
    ff_ram[9035] = 8'h00;
    ff_ram[9036] = 8'h00;
    ff_ram[9037] = 8'h00;
    ff_ram[9038] = 8'h00;
    ff_ram[9039] = 8'h00;
    ff_ram[9040] = 8'h00;
    ff_ram[9041] = 8'h00;
    ff_ram[9042] = 8'h00;
    ff_ram[9043] = 8'h00;
    ff_ram[9044] = 8'h00;
    ff_ram[9045] = 8'h00;
    ff_ram[9046] = 8'h00;
    ff_ram[9047] = 8'h00;
    ff_ram[9048] = 8'h00;
    ff_ram[9049] = 8'h00;
    ff_ram[9050] = 8'h00;
    ff_ram[9051] = 8'h00;
    ff_ram[9052] = 8'h00;
    ff_ram[9053] = 8'h00;
    ff_ram[9054] = 8'h00;
    ff_ram[9055] = 8'h00;
    ff_ram[9056] = 8'h00;
    ff_ram[9057] = 8'h00;
    ff_ram[9058] = 8'h00;
    ff_ram[9059] = 8'h00;
    ff_ram[9060] = 8'h00;
    ff_ram[9061] = 8'h00;
    ff_ram[9062] = 8'h00;
    ff_ram[9063] = 8'h00;
    ff_ram[9064] = 8'h00;
    ff_ram[9065] = 8'h00;
    ff_ram[9066] = 8'h00;
    ff_ram[9067] = 8'h00;
    ff_ram[9068] = 8'h00;
    ff_ram[9069] = 8'h00;
    ff_ram[9070] = 8'h00;
    ff_ram[9071] = 8'h00;
    ff_ram[9072] = 8'h00;
    ff_ram[9073] = 8'h00;
    ff_ram[9074] = 8'h00;
    ff_ram[9075] = 8'h00;
    ff_ram[9076] = 8'h00;
    ff_ram[9077] = 8'h00;
    ff_ram[9078] = 8'h00;
    ff_ram[9079] = 8'h00;
    ff_ram[9080] = 8'h00;
    ff_ram[9081] = 8'h00;
    ff_ram[9082] = 8'h00;
    ff_ram[9083] = 8'h00;
    ff_ram[9084] = 8'h00;
    ff_ram[9085] = 8'h00;
    ff_ram[9086] = 8'h00;
    ff_ram[9087] = 8'h00;
    ff_ram[9088] = 8'h00;
    ff_ram[9089] = 8'h00;
    ff_ram[9090] = 8'h00;
    ff_ram[9091] = 8'h00;
    ff_ram[9092] = 8'h00;
    ff_ram[9093] = 8'h00;
    ff_ram[9094] = 8'h00;
    ff_ram[9095] = 8'h00;
    ff_ram[9096] = 8'h00;
    ff_ram[9097] = 8'h00;
    ff_ram[9098] = 8'h00;
    ff_ram[9099] = 8'h00;
    ff_ram[9100] = 8'h00;
    ff_ram[9101] = 8'h00;
    ff_ram[9102] = 8'h00;
    ff_ram[9103] = 8'h00;
    ff_ram[9104] = 8'h00;
    ff_ram[9105] = 8'h00;
    ff_ram[9106] = 8'h00;
    ff_ram[9107] = 8'h00;
    ff_ram[9108] = 8'h00;
    ff_ram[9109] = 8'h00;
    ff_ram[9110] = 8'h00;
    ff_ram[9111] = 8'h00;
    ff_ram[9112] = 8'h00;
    ff_ram[9113] = 8'h00;
    ff_ram[9114] = 8'h00;
    ff_ram[9115] = 8'h00;
    ff_ram[9116] = 8'h00;
    ff_ram[9117] = 8'h00;
    ff_ram[9118] = 8'h00;
    ff_ram[9119] = 8'h00;
    ff_ram[9120] = 8'h00;
    ff_ram[9121] = 8'h00;
    ff_ram[9122] = 8'h00;
    ff_ram[9123] = 8'h00;
    ff_ram[9124] = 8'h00;
    ff_ram[9125] = 8'h00;
    ff_ram[9126] = 8'h00;
    ff_ram[9127] = 8'h00;
    ff_ram[9128] = 8'h00;
    ff_ram[9129] = 8'h00;
    ff_ram[9130] = 8'h00;
    ff_ram[9131] = 8'h00;
    ff_ram[9132] = 8'h00;
    ff_ram[9133] = 8'h00;
    ff_ram[9134] = 8'h00;
    ff_ram[9135] = 8'h00;
    ff_ram[9136] = 8'h00;
    ff_ram[9137] = 8'h00;
    ff_ram[9138] = 8'h00;
    ff_ram[9139] = 8'h00;
    ff_ram[9140] = 8'h00;
    ff_ram[9141] = 8'h00;
    ff_ram[9142] = 8'h00;
    ff_ram[9143] = 8'h00;
    ff_ram[9144] = 8'h00;
    ff_ram[9145] = 8'h00;
    ff_ram[9146] = 8'h00;
    ff_ram[9147] = 8'h00;
    ff_ram[9148] = 8'h00;
    ff_ram[9149] = 8'h00;
    ff_ram[9150] = 8'h00;
    ff_ram[9151] = 8'h00;
    ff_ram[9152] = 8'h00;
    ff_ram[9153] = 8'h00;
    ff_ram[9154] = 8'h00;
    ff_ram[9155] = 8'h00;
    ff_ram[9156] = 8'h00;
    ff_ram[9157] = 8'h00;
    ff_ram[9158] = 8'h00;
    ff_ram[9159] = 8'h00;
    ff_ram[9160] = 8'h00;
    ff_ram[9161] = 8'h00;
    ff_ram[9162] = 8'h00;
    ff_ram[9163] = 8'h00;
    ff_ram[9164] = 8'h00;
    ff_ram[9165] = 8'h00;
    ff_ram[9166] = 8'h00;
    ff_ram[9167] = 8'h00;
    ff_ram[9168] = 8'h00;
    ff_ram[9169] = 8'h00;
    ff_ram[9170] = 8'h00;
    ff_ram[9171] = 8'h00;
    ff_ram[9172] = 8'h00;
    ff_ram[9173] = 8'h00;
    ff_ram[9174] = 8'h00;
    ff_ram[9175] = 8'h00;
    ff_ram[9176] = 8'h00;
    ff_ram[9177] = 8'h00;
    ff_ram[9178] = 8'h00;
    ff_ram[9179] = 8'h00;
    ff_ram[9180] = 8'h00;
    ff_ram[9181] = 8'h00;
    ff_ram[9182] = 8'h00;
    ff_ram[9183] = 8'h00;
    ff_ram[9184] = 8'h00;
    ff_ram[9185] = 8'h00;
    ff_ram[9186] = 8'h00;
    ff_ram[9187] = 8'h00;
    ff_ram[9188] = 8'h00;
    ff_ram[9189] = 8'h00;
    ff_ram[9190] = 8'h00;
    ff_ram[9191] = 8'h00;
    ff_ram[9192] = 8'h00;
    ff_ram[9193] = 8'h00;
    ff_ram[9194] = 8'h00;
    ff_ram[9195] = 8'h00;
    ff_ram[9196] = 8'h00;
    ff_ram[9197] = 8'h00;
    ff_ram[9198] = 8'h00;
    ff_ram[9199] = 8'h00;
    ff_ram[9200] = 8'h00;
    ff_ram[9201] = 8'h00;
    ff_ram[9202] = 8'h00;
    ff_ram[9203] = 8'h00;
    ff_ram[9204] = 8'h00;
    ff_ram[9205] = 8'h00;
    ff_ram[9206] = 8'h00;
    ff_ram[9207] = 8'h00;
    ff_ram[9208] = 8'h00;
    ff_ram[9209] = 8'h00;
    ff_ram[9210] = 8'h00;
    ff_ram[9211] = 8'h00;
    ff_ram[9212] = 8'h00;
    ff_ram[9213] = 8'h00;
    ff_ram[9214] = 8'h00;
    ff_ram[9215] = 8'h00;
    ff_ram[9216] = 8'h00;
    ff_ram[9217] = 8'h00;
    ff_ram[9218] = 8'h00;
    ff_ram[9219] = 8'h00;
    ff_ram[9220] = 8'h00;
    ff_ram[9221] = 8'h00;
    ff_ram[9222] = 8'h00;
    ff_ram[9223] = 8'h00;
    ff_ram[9224] = 8'h00;
    ff_ram[9225] = 8'h00;
    ff_ram[9226] = 8'h00;
    ff_ram[9227] = 8'h00;
    ff_ram[9228] = 8'h00;
    ff_ram[9229] = 8'h00;
    ff_ram[9230] = 8'h00;
    ff_ram[9231] = 8'h00;
    ff_ram[9232] = 8'h00;
    ff_ram[9233] = 8'h00;
    ff_ram[9234] = 8'h00;
    ff_ram[9235] = 8'h00;
    ff_ram[9236] = 8'h00;
    ff_ram[9237] = 8'h00;
    ff_ram[9238] = 8'h00;
    ff_ram[9239] = 8'h00;
    ff_ram[9240] = 8'h00;
    ff_ram[9241] = 8'h00;
    ff_ram[9242] = 8'h00;
    ff_ram[9243] = 8'h00;
    ff_ram[9244] = 8'h00;
    ff_ram[9245] = 8'h00;
    ff_ram[9246] = 8'h00;
    ff_ram[9247] = 8'h00;
    ff_ram[9248] = 8'h00;
    ff_ram[9249] = 8'h00;
    ff_ram[9250] = 8'h00;
    ff_ram[9251] = 8'h00;
    ff_ram[9252] = 8'h00;
    ff_ram[9253] = 8'h00;
    ff_ram[9254] = 8'h00;
    ff_ram[9255] = 8'h00;
    ff_ram[9256] = 8'h00;
    ff_ram[9257] = 8'h00;
    ff_ram[9258] = 8'h00;
    ff_ram[9259] = 8'h00;
    ff_ram[9260] = 8'h00;
    ff_ram[9261] = 8'h00;
    ff_ram[9262] = 8'h00;
    ff_ram[9263] = 8'h00;
    ff_ram[9264] = 8'h00;
    ff_ram[9265] = 8'h00;
    ff_ram[9266] = 8'h00;
    ff_ram[9267] = 8'h00;
    ff_ram[9268] = 8'h00;
    ff_ram[9269] = 8'h00;
    ff_ram[9270] = 8'h00;
    ff_ram[9271] = 8'h00;
    ff_ram[9272] = 8'h00;
    ff_ram[9273] = 8'h00;
    ff_ram[9274] = 8'h00;
    ff_ram[9275] = 8'h00;
    ff_ram[9276] = 8'h00;
    ff_ram[9277] = 8'h00;
    ff_ram[9278] = 8'h00;
    ff_ram[9279] = 8'h00;
    ff_ram[9280] = 8'h00;
    ff_ram[9281] = 8'h00;
    ff_ram[9282] = 8'h00;
    ff_ram[9283] = 8'h00;
    ff_ram[9284] = 8'h00;
    ff_ram[9285] = 8'h00;
    ff_ram[9286] = 8'h00;
    ff_ram[9287] = 8'h00;
    ff_ram[9288] = 8'h00;
    ff_ram[9289] = 8'h00;
    ff_ram[9290] = 8'h00;
    ff_ram[9291] = 8'h00;
    ff_ram[9292] = 8'h00;
    ff_ram[9293] = 8'h00;
    ff_ram[9294] = 8'h00;
    ff_ram[9295] = 8'h00;
    ff_ram[9296] = 8'h00;
    ff_ram[9297] = 8'h00;
    ff_ram[9298] = 8'h00;
    ff_ram[9299] = 8'h00;
    ff_ram[9300] = 8'h00;
    ff_ram[9301] = 8'h00;
    ff_ram[9302] = 8'h00;
    ff_ram[9303] = 8'h00;
    ff_ram[9304] = 8'h00;
    ff_ram[9305] = 8'h00;
    ff_ram[9306] = 8'h00;
    ff_ram[9307] = 8'h00;
    ff_ram[9308] = 8'h00;
    ff_ram[9309] = 8'h00;
    ff_ram[9310] = 8'h00;
    ff_ram[9311] = 8'h00;
    ff_ram[9312] = 8'h00;
    ff_ram[9313] = 8'h00;
    ff_ram[9314] = 8'h00;
    ff_ram[9315] = 8'h00;
    ff_ram[9316] = 8'h00;
    ff_ram[9317] = 8'h00;
    ff_ram[9318] = 8'h00;
    ff_ram[9319] = 8'h00;
    ff_ram[9320] = 8'h00;
    ff_ram[9321] = 8'h00;
    ff_ram[9322] = 8'h00;
    ff_ram[9323] = 8'h00;
    ff_ram[9324] = 8'h00;
    ff_ram[9325] = 8'h00;
    ff_ram[9326] = 8'h00;
    ff_ram[9327] = 8'h00;
    ff_ram[9328] = 8'h00;
    ff_ram[9329] = 8'h00;
    ff_ram[9330] = 8'h00;
    ff_ram[9331] = 8'h00;
    ff_ram[9332] = 8'h00;
    ff_ram[9333] = 8'h00;
    ff_ram[9334] = 8'h00;
    ff_ram[9335] = 8'h00;
    ff_ram[9336] = 8'h00;
    ff_ram[9337] = 8'h00;
    ff_ram[9338] = 8'h00;
    ff_ram[9339] = 8'h00;
    ff_ram[9340] = 8'h00;
    ff_ram[9341] = 8'h00;
    ff_ram[9342] = 8'h00;
    ff_ram[9343] = 8'h00;
    ff_ram[9344] = 8'h00;
    ff_ram[9345] = 8'h00;
    ff_ram[9346] = 8'h00;
    ff_ram[9347] = 8'h00;
    ff_ram[9348] = 8'h00;
    ff_ram[9349] = 8'h00;
    ff_ram[9350] = 8'h00;
    ff_ram[9351] = 8'h00;
    ff_ram[9352] = 8'h00;
    ff_ram[9353] = 8'h00;
    ff_ram[9354] = 8'h00;
    ff_ram[9355] = 8'h00;
    ff_ram[9356] = 8'h00;
    ff_ram[9357] = 8'h00;
    ff_ram[9358] = 8'h00;
    ff_ram[9359] = 8'h00;
    ff_ram[9360] = 8'h00;
    ff_ram[9361] = 8'h00;
    ff_ram[9362] = 8'h00;
    ff_ram[9363] = 8'h00;
    ff_ram[9364] = 8'h00;
    ff_ram[9365] = 8'h00;
    ff_ram[9366] = 8'h00;
    ff_ram[9367] = 8'h00;
    ff_ram[9368] = 8'h00;
    ff_ram[9369] = 8'h00;
    ff_ram[9370] = 8'h00;
    ff_ram[9371] = 8'h00;
    ff_ram[9372] = 8'h00;
    ff_ram[9373] = 8'h00;
    ff_ram[9374] = 8'h00;
    ff_ram[9375] = 8'h00;
    ff_ram[9376] = 8'h00;
    ff_ram[9377] = 8'h00;
    ff_ram[9378] = 8'h00;
    ff_ram[9379] = 8'h00;
    ff_ram[9380] = 8'h00;
    ff_ram[9381] = 8'h00;
    ff_ram[9382] = 8'h00;
    ff_ram[9383] = 8'h00;
    ff_ram[9384] = 8'h00;
    ff_ram[9385] = 8'h00;
    ff_ram[9386] = 8'h00;
    ff_ram[9387] = 8'h00;
    ff_ram[9388] = 8'h00;
    ff_ram[9389] = 8'h00;
    ff_ram[9390] = 8'h00;
    ff_ram[9391] = 8'h00;
    ff_ram[9392] = 8'h00;
    ff_ram[9393] = 8'h00;
    ff_ram[9394] = 8'h00;
    ff_ram[9395] = 8'h00;
    ff_ram[9396] = 8'h00;
    ff_ram[9397] = 8'h00;
    ff_ram[9398] = 8'h00;
    ff_ram[9399] = 8'h00;
    ff_ram[9400] = 8'h00;
    ff_ram[9401] = 8'h00;
    ff_ram[9402] = 8'h00;
    ff_ram[9403] = 8'h00;
    ff_ram[9404] = 8'h00;
    ff_ram[9405] = 8'h00;
    ff_ram[9406] = 8'h00;
    ff_ram[9407] = 8'h00;
    ff_ram[9408] = 8'h00;
    ff_ram[9409] = 8'h00;
    ff_ram[9410] = 8'h00;
    ff_ram[9411] = 8'h00;
    ff_ram[9412] = 8'h00;
    ff_ram[9413] = 8'h00;
    ff_ram[9414] = 8'h00;
    ff_ram[9415] = 8'h00;
    ff_ram[9416] = 8'h00;
    ff_ram[9417] = 8'h00;
    ff_ram[9418] = 8'h00;
    ff_ram[9419] = 8'h00;
    ff_ram[9420] = 8'h00;
    ff_ram[9421] = 8'h00;
    ff_ram[9422] = 8'h00;
    ff_ram[9423] = 8'h00;
    ff_ram[9424] = 8'h00;
    ff_ram[9425] = 8'h00;
    ff_ram[9426] = 8'h00;
    ff_ram[9427] = 8'h00;
    ff_ram[9428] = 8'h00;
    ff_ram[9429] = 8'h00;
    ff_ram[9430] = 8'h00;
    ff_ram[9431] = 8'h00;
    ff_ram[9432] = 8'h00;
    ff_ram[9433] = 8'h00;
    ff_ram[9434] = 8'h00;
    ff_ram[9435] = 8'h00;
    ff_ram[9436] = 8'h00;
    ff_ram[9437] = 8'h00;
    ff_ram[9438] = 8'h00;
    ff_ram[9439] = 8'h00;
    ff_ram[9440] = 8'h00;
    ff_ram[9441] = 8'h00;
    ff_ram[9442] = 8'h00;
    ff_ram[9443] = 8'h00;
    ff_ram[9444] = 8'h00;
    ff_ram[9445] = 8'h00;
    ff_ram[9446] = 8'h00;
    ff_ram[9447] = 8'h00;
    ff_ram[9448] = 8'h00;
    ff_ram[9449] = 8'h00;
    ff_ram[9450] = 8'h00;
    ff_ram[9451] = 8'h00;
    ff_ram[9452] = 8'h00;
    ff_ram[9453] = 8'h00;
    ff_ram[9454] = 8'h00;
    ff_ram[9455] = 8'h00;
    ff_ram[9456] = 8'h00;
    ff_ram[9457] = 8'h00;
    ff_ram[9458] = 8'h00;
    ff_ram[9459] = 8'h00;
    ff_ram[9460] = 8'h00;
    ff_ram[9461] = 8'h00;
    ff_ram[9462] = 8'h00;
    ff_ram[9463] = 8'h00;
    ff_ram[9464] = 8'h00;
    ff_ram[9465] = 8'h00;
    ff_ram[9466] = 8'h00;
    ff_ram[9467] = 8'h00;
    ff_ram[9468] = 8'h00;
    ff_ram[9469] = 8'h00;
    ff_ram[9470] = 8'h00;
    ff_ram[9471] = 8'h00;
    ff_ram[9472] = 8'h00;
    ff_ram[9473] = 8'h00;
    ff_ram[9474] = 8'h00;
    ff_ram[9475] = 8'h00;
    ff_ram[9476] = 8'h00;
    ff_ram[9477] = 8'h00;
    ff_ram[9478] = 8'h00;
    ff_ram[9479] = 8'h00;
    ff_ram[9480] = 8'h00;
    ff_ram[9481] = 8'h00;
    ff_ram[9482] = 8'h00;
    ff_ram[9483] = 8'h00;
    ff_ram[9484] = 8'h00;
    ff_ram[9485] = 8'h00;
    ff_ram[9486] = 8'h00;
    ff_ram[9487] = 8'h00;
    ff_ram[9488] = 8'h00;
    ff_ram[9489] = 8'h00;
    ff_ram[9490] = 8'h00;
    ff_ram[9491] = 8'h00;
    ff_ram[9492] = 8'h00;
    ff_ram[9493] = 8'h00;
    ff_ram[9494] = 8'h00;
    ff_ram[9495] = 8'h00;
    ff_ram[9496] = 8'h00;
    ff_ram[9497] = 8'h00;
    ff_ram[9498] = 8'h00;
    ff_ram[9499] = 8'h00;
    ff_ram[9500] = 8'h00;
    ff_ram[9501] = 8'h00;
    ff_ram[9502] = 8'h00;
    ff_ram[9503] = 8'h00;
    ff_ram[9504] = 8'h00;
    ff_ram[9505] = 8'h00;
    ff_ram[9506] = 8'h00;
    ff_ram[9507] = 8'h00;
    ff_ram[9508] = 8'h00;
    ff_ram[9509] = 8'h00;
    ff_ram[9510] = 8'h00;
    ff_ram[9511] = 8'h00;
    ff_ram[9512] = 8'h00;
    ff_ram[9513] = 8'h00;
    ff_ram[9514] = 8'h00;
    ff_ram[9515] = 8'h00;
    ff_ram[9516] = 8'h00;
    ff_ram[9517] = 8'h00;
    ff_ram[9518] = 8'h00;
    ff_ram[9519] = 8'h00;
    ff_ram[9520] = 8'h00;
    ff_ram[9521] = 8'h00;
    ff_ram[9522] = 8'h00;
    ff_ram[9523] = 8'h00;
    ff_ram[9524] = 8'h00;
    ff_ram[9525] = 8'h00;
    ff_ram[9526] = 8'h00;
    ff_ram[9527] = 8'h00;
    ff_ram[9528] = 8'h00;
    ff_ram[9529] = 8'h00;
    ff_ram[9530] = 8'h00;
    ff_ram[9531] = 8'h00;
    ff_ram[9532] = 8'h00;
    ff_ram[9533] = 8'h00;
    ff_ram[9534] = 8'h00;
    ff_ram[9535] = 8'h00;
    ff_ram[9536] = 8'h00;
    ff_ram[9537] = 8'h00;
    ff_ram[9538] = 8'h00;
    ff_ram[9539] = 8'h00;
    ff_ram[9540] = 8'h00;
    ff_ram[9541] = 8'h00;
    ff_ram[9542] = 8'h00;
    ff_ram[9543] = 8'h00;
    ff_ram[9544] = 8'h00;
    ff_ram[9545] = 8'h00;
    ff_ram[9546] = 8'h00;
    ff_ram[9547] = 8'h00;
    ff_ram[9548] = 8'h00;
    ff_ram[9549] = 8'h00;
    ff_ram[9550] = 8'h00;
    ff_ram[9551] = 8'h00;
    ff_ram[9552] = 8'h00;
    ff_ram[9553] = 8'h00;
    ff_ram[9554] = 8'h00;
    ff_ram[9555] = 8'h00;
    ff_ram[9556] = 8'h00;
    ff_ram[9557] = 8'h00;
    ff_ram[9558] = 8'h00;
    ff_ram[9559] = 8'h00;
    ff_ram[9560] = 8'h00;
    ff_ram[9561] = 8'h00;
    ff_ram[9562] = 8'h00;
    ff_ram[9563] = 8'h00;
    ff_ram[9564] = 8'h00;
    ff_ram[9565] = 8'h00;
    ff_ram[9566] = 8'h00;
    ff_ram[9567] = 8'h00;
    ff_ram[9568] = 8'h00;
    ff_ram[9569] = 8'h00;
    ff_ram[9570] = 8'h00;
    ff_ram[9571] = 8'h00;
    ff_ram[9572] = 8'h00;
    ff_ram[9573] = 8'h00;
    ff_ram[9574] = 8'h00;
    ff_ram[9575] = 8'h00;
    ff_ram[9576] = 8'h00;
    ff_ram[9577] = 8'h00;
    ff_ram[9578] = 8'h00;
    ff_ram[9579] = 8'h00;
    ff_ram[9580] = 8'h00;
    ff_ram[9581] = 8'h00;
    ff_ram[9582] = 8'h00;
    ff_ram[9583] = 8'h00;
    ff_ram[9584] = 8'h00;
    ff_ram[9585] = 8'h00;
    ff_ram[9586] = 8'h00;
    ff_ram[9587] = 8'h00;
    ff_ram[9588] = 8'h00;
    ff_ram[9589] = 8'h00;
    ff_ram[9590] = 8'h00;
    ff_ram[9591] = 8'h00;
    ff_ram[9592] = 8'h00;
    ff_ram[9593] = 8'h00;
    ff_ram[9594] = 8'h00;
    ff_ram[9595] = 8'h00;
    ff_ram[9596] = 8'h00;
    ff_ram[9597] = 8'h00;
    ff_ram[9598] = 8'h00;
    ff_ram[9599] = 8'h00;
    ff_ram[9600] = 8'h00;
    ff_ram[9601] = 8'h00;
    ff_ram[9602] = 8'h00;
    ff_ram[9603] = 8'h00;
    ff_ram[9604] = 8'h00;
    ff_ram[9605] = 8'h00;
    ff_ram[9606] = 8'h00;
    ff_ram[9607] = 8'h00;
    ff_ram[9608] = 8'h00;
    ff_ram[9609] = 8'h00;
    ff_ram[9610] = 8'h00;
    ff_ram[9611] = 8'h00;
    ff_ram[9612] = 8'h00;
    ff_ram[9613] = 8'h00;
    ff_ram[9614] = 8'h00;
    ff_ram[9615] = 8'h00;
    ff_ram[9616] = 8'h00;
    ff_ram[9617] = 8'h00;
    ff_ram[9618] = 8'h00;
    ff_ram[9619] = 8'h00;
    ff_ram[9620] = 8'h00;
    ff_ram[9621] = 8'h00;
    ff_ram[9622] = 8'h00;
    ff_ram[9623] = 8'h00;
    ff_ram[9624] = 8'h00;
    ff_ram[9625] = 8'h00;
    ff_ram[9626] = 8'h00;
    ff_ram[9627] = 8'h00;
    ff_ram[9628] = 8'h00;
    ff_ram[9629] = 8'h00;
    ff_ram[9630] = 8'h00;
    ff_ram[9631] = 8'h00;
    ff_ram[9632] = 8'h00;
    ff_ram[9633] = 8'h00;
    ff_ram[9634] = 8'h00;
    ff_ram[9635] = 8'h00;
    ff_ram[9636] = 8'h00;
    ff_ram[9637] = 8'h00;
    ff_ram[9638] = 8'h00;
    ff_ram[9639] = 8'h00;
    ff_ram[9640] = 8'h00;
    ff_ram[9641] = 8'h00;
    ff_ram[9642] = 8'h00;
    ff_ram[9643] = 8'h00;
    ff_ram[9644] = 8'h00;
    ff_ram[9645] = 8'h00;
    ff_ram[9646] = 8'h00;
    ff_ram[9647] = 8'h00;
    ff_ram[9648] = 8'h00;
    ff_ram[9649] = 8'h00;
    ff_ram[9650] = 8'h00;
    ff_ram[9651] = 8'h00;
    ff_ram[9652] = 8'h00;
    ff_ram[9653] = 8'h00;
    ff_ram[9654] = 8'h00;
    ff_ram[9655] = 8'h00;
    ff_ram[9656] = 8'h00;
    ff_ram[9657] = 8'h00;
    ff_ram[9658] = 8'h00;
    ff_ram[9659] = 8'h00;
    ff_ram[9660] = 8'h00;
    ff_ram[9661] = 8'h00;
    ff_ram[9662] = 8'h00;
    ff_ram[9663] = 8'h00;
    ff_ram[9664] = 8'h00;
    ff_ram[9665] = 8'h00;
    ff_ram[9666] = 8'h00;
    ff_ram[9667] = 8'h00;
    ff_ram[9668] = 8'h00;
    ff_ram[9669] = 8'h00;
    ff_ram[9670] = 8'h00;
    ff_ram[9671] = 8'h00;
    ff_ram[9672] = 8'h00;
    ff_ram[9673] = 8'h00;
    ff_ram[9674] = 8'h00;
    ff_ram[9675] = 8'h00;
    ff_ram[9676] = 8'h00;
    ff_ram[9677] = 8'h00;
    ff_ram[9678] = 8'h00;
    ff_ram[9679] = 8'h00;
    ff_ram[9680] = 8'h00;
    ff_ram[9681] = 8'h00;
    ff_ram[9682] = 8'h00;
    ff_ram[9683] = 8'h00;
    ff_ram[9684] = 8'h00;
    ff_ram[9685] = 8'h00;
    ff_ram[9686] = 8'h00;
    ff_ram[9687] = 8'h00;
    ff_ram[9688] = 8'h00;
    ff_ram[9689] = 8'h00;
    ff_ram[9690] = 8'h00;
    ff_ram[9691] = 8'h00;
    ff_ram[9692] = 8'h00;
    ff_ram[9693] = 8'h00;
    ff_ram[9694] = 8'h00;
    ff_ram[9695] = 8'h00;
    ff_ram[9696] = 8'h00;
    ff_ram[9697] = 8'h00;
    ff_ram[9698] = 8'h00;
    ff_ram[9699] = 8'h00;
    ff_ram[9700] = 8'h00;
    ff_ram[9701] = 8'h00;
    ff_ram[9702] = 8'h00;
    ff_ram[9703] = 8'h00;
    ff_ram[9704] = 8'h00;
    ff_ram[9705] = 8'h00;
    ff_ram[9706] = 8'h00;
    ff_ram[9707] = 8'h00;
    ff_ram[9708] = 8'h00;
    ff_ram[9709] = 8'h00;
    ff_ram[9710] = 8'h00;
    ff_ram[9711] = 8'h00;
    ff_ram[9712] = 8'h00;
    ff_ram[9713] = 8'h00;
    ff_ram[9714] = 8'h00;
    ff_ram[9715] = 8'h00;
    ff_ram[9716] = 8'h00;
    ff_ram[9717] = 8'h00;
    ff_ram[9718] = 8'h00;
    ff_ram[9719] = 8'h00;
    ff_ram[9720] = 8'h00;
    ff_ram[9721] = 8'h00;
    ff_ram[9722] = 8'h00;
    ff_ram[9723] = 8'h00;
    ff_ram[9724] = 8'h00;
    ff_ram[9725] = 8'h00;
    ff_ram[9726] = 8'h00;
    ff_ram[9727] = 8'h00;
    ff_ram[9728] = 8'h00;
    ff_ram[9729] = 8'h00;
    ff_ram[9730] = 8'h00;
    ff_ram[9731] = 8'h00;
    ff_ram[9732] = 8'h00;
    ff_ram[9733] = 8'h00;
    ff_ram[9734] = 8'h00;
    ff_ram[9735] = 8'h00;
    ff_ram[9736] = 8'h00;
    ff_ram[9737] = 8'h00;
    ff_ram[9738] = 8'h00;
    ff_ram[9739] = 8'h00;
    ff_ram[9740] = 8'h00;
    ff_ram[9741] = 8'h00;
    ff_ram[9742] = 8'h00;
    ff_ram[9743] = 8'h00;
    ff_ram[9744] = 8'h00;
    ff_ram[9745] = 8'h00;
    ff_ram[9746] = 8'h00;
    ff_ram[9747] = 8'h00;
    ff_ram[9748] = 8'h00;
    ff_ram[9749] = 8'h00;
    ff_ram[9750] = 8'h00;
    ff_ram[9751] = 8'h00;
    ff_ram[9752] = 8'h00;
    ff_ram[9753] = 8'h00;
    ff_ram[9754] = 8'h00;
    ff_ram[9755] = 8'h00;
    ff_ram[9756] = 8'h00;
    ff_ram[9757] = 8'h00;
    ff_ram[9758] = 8'h00;
    ff_ram[9759] = 8'h00;
    ff_ram[9760] = 8'h00;
    ff_ram[9761] = 8'h00;
    ff_ram[9762] = 8'h00;
    ff_ram[9763] = 8'h00;
    ff_ram[9764] = 8'h00;
    ff_ram[9765] = 8'h00;
    ff_ram[9766] = 8'h00;
    ff_ram[9767] = 8'h00;
    ff_ram[9768] = 8'h00;
    ff_ram[9769] = 8'h00;
    ff_ram[9770] = 8'h00;
    ff_ram[9771] = 8'h00;
    ff_ram[9772] = 8'h00;
    ff_ram[9773] = 8'h00;
    ff_ram[9774] = 8'h00;
    ff_ram[9775] = 8'h00;
    ff_ram[9776] = 8'h00;
    ff_ram[9777] = 8'h00;
    ff_ram[9778] = 8'h00;
    ff_ram[9779] = 8'h00;
    ff_ram[9780] = 8'h00;
    ff_ram[9781] = 8'h00;
    ff_ram[9782] = 8'h00;
    ff_ram[9783] = 8'h00;
    ff_ram[9784] = 8'h00;
    ff_ram[9785] = 8'h00;
    ff_ram[9786] = 8'h00;
    ff_ram[9787] = 8'h00;
    ff_ram[9788] = 8'h00;
    ff_ram[9789] = 8'h00;
    ff_ram[9790] = 8'h00;
    ff_ram[9791] = 8'h00;
    ff_ram[9792] = 8'h00;
    ff_ram[9793] = 8'h00;
    ff_ram[9794] = 8'h00;
    ff_ram[9795] = 8'h00;
    ff_ram[9796] = 8'h00;
    ff_ram[9797] = 8'h00;
    ff_ram[9798] = 8'h00;
    ff_ram[9799] = 8'h00;
    ff_ram[9800] = 8'h00;
    ff_ram[9801] = 8'h00;
    ff_ram[9802] = 8'h00;
    ff_ram[9803] = 8'h00;
    ff_ram[9804] = 8'h00;
    ff_ram[9805] = 8'h00;
    ff_ram[9806] = 8'h00;
    ff_ram[9807] = 8'h00;
    ff_ram[9808] = 8'h00;
    ff_ram[9809] = 8'h00;
    ff_ram[9810] = 8'h00;
    ff_ram[9811] = 8'h00;
    ff_ram[9812] = 8'h00;
    ff_ram[9813] = 8'h00;
    ff_ram[9814] = 8'h00;
    ff_ram[9815] = 8'h00;
    ff_ram[9816] = 8'h00;
    ff_ram[9817] = 8'h00;
    ff_ram[9818] = 8'h00;
    ff_ram[9819] = 8'h00;
    ff_ram[9820] = 8'h00;
    ff_ram[9821] = 8'h00;
    ff_ram[9822] = 8'h00;
    ff_ram[9823] = 8'h00;
    ff_ram[9824] = 8'h00;
    ff_ram[9825] = 8'h00;
    ff_ram[9826] = 8'h00;
    ff_ram[9827] = 8'h00;
    ff_ram[9828] = 8'h00;
    ff_ram[9829] = 8'h00;
    ff_ram[9830] = 8'h00;
    ff_ram[9831] = 8'h00;
    ff_ram[9832] = 8'h00;
    ff_ram[9833] = 8'h00;
    ff_ram[9834] = 8'h00;
    ff_ram[9835] = 8'h00;
    ff_ram[9836] = 8'h00;
    ff_ram[9837] = 8'h00;
    ff_ram[9838] = 8'h00;
    ff_ram[9839] = 8'h00;
    ff_ram[9840] = 8'h00;
    ff_ram[9841] = 8'h00;
    ff_ram[9842] = 8'h00;
    ff_ram[9843] = 8'h00;
    ff_ram[9844] = 8'h00;
    ff_ram[9845] = 8'h00;
    ff_ram[9846] = 8'h00;
    ff_ram[9847] = 8'h00;
    ff_ram[9848] = 8'h00;
    ff_ram[9849] = 8'h00;
    ff_ram[9850] = 8'h00;
    ff_ram[9851] = 8'h00;
    ff_ram[9852] = 8'h00;
    ff_ram[9853] = 8'h00;
    ff_ram[9854] = 8'h00;
    ff_ram[9855] = 8'h00;
    ff_ram[9856] = 8'h00;
    ff_ram[9857] = 8'h00;
    ff_ram[9858] = 8'h00;
    ff_ram[9859] = 8'h00;
    ff_ram[9860] = 8'h00;
    ff_ram[9861] = 8'h00;
    ff_ram[9862] = 8'h00;
    ff_ram[9863] = 8'h00;
    ff_ram[9864] = 8'h00;
    ff_ram[9865] = 8'h00;
    ff_ram[9866] = 8'h00;
    ff_ram[9867] = 8'h00;
    ff_ram[9868] = 8'h00;
    ff_ram[9869] = 8'h00;
    ff_ram[9870] = 8'h00;
    ff_ram[9871] = 8'h00;
    ff_ram[9872] = 8'h00;
    ff_ram[9873] = 8'h00;
    ff_ram[9874] = 8'h00;
    ff_ram[9875] = 8'h00;
    ff_ram[9876] = 8'h00;
    ff_ram[9877] = 8'h00;
    ff_ram[9878] = 8'h00;
    ff_ram[9879] = 8'h00;
    ff_ram[9880] = 8'h00;
    ff_ram[9881] = 8'h00;
    ff_ram[9882] = 8'h00;
    ff_ram[9883] = 8'h00;
    ff_ram[9884] = 8'h00;
    ff_ram[9885] = 8'h00;
    ff_ram[9886] = 8'h00;
    ff_ram[9887] = 8'h00;
    ff_ram[9888] = 8'h00;
    ff_ram[9889] = 8'h00;
    ff_ram[9890] = 8'h00;
    ff_ram[9891] = 8'h00;
    ff_ram[9892] = 8'h00;
    ff_ram[9893] = 8'h00;
    ff_ram[9894] = 8'h00;
    ff_ram[9895] = 8'h00;
    ff_ram[9896] = 8'h00;
    ff_ram[9897] = 8'h00;
    ff_ram[9898] = 8'h00;
    ff_ram[9899] = 8'h00;
    ff_ram[9900] = 8'h00;
    ff_ram[9901] = 8'h00;
    ff_ram[9902] = 8'h00;
    ff_ram[9903] = 8'h00;
    ff_ram[9904] = 8'h00;
    ff_ram[9905] = 8'h00;
    ff_ram[9906] = 8'h00;
    ff_ram[9907] = 8'h00;
    ff_ram[9908] = 8'h00;
    ff_ram[9909] = 8'h00;
    ff_ram[9910] = 8'h00;
    ff_ram[9911] = 8'h00;
    ff_ram[9912] = 8'h00;
    ff_ram[9913] = 8'h00;
    ff_ram[9914] = 8'h00;
    ff_ram[9915] = 8'h00;
    ff_ram[9916] = 8'h00;
    ff_ram[9917] = 8'h00;
    ff_ram[9918] = 8'h00;
    ff_ram[9919] = 8'h00;
    ff_ram[9920] = 8'h00;
    ff_ram[9921] = 8'h00;
    ff_ram[9922] = 8'h00;
    ff_ram[9923] = 8'h00;
    ff_ram[9924] = 8'h00;
    ff_ram[9925] = 8'h00;
    ff_ram[9926] = 8'h00;
    ff_ram[9927] = 8'h00;
    ff_ram[9928] = 8'h00;
    ff_ram[9929] = 8'h00;
    ff_ram[9930] = 8'h00;
    ff_ram[9931] = 8'h00;
    ff_ram[9932] = 8'h00;
    ff_ram[9933] = 8'h00;
    ff_ram[9934] = 8'h00;
    ff_ram[9935] = 8'h00;
    ff_ram[9936] = 8'h00;
    ff_ram[9937] = 8'h00;
    ff_ram[9938] = 8'h00;
    ff_ram[9939] = 8'h00;
    ff_ram[9940] = 8'h00;
    ff_ram[9941] = 8'h00;
    ff_ram[9942] = 8'h00;
    ff_ram[9943] = 8'h00;
    ff_ram[9944] = 8'h00;
    ff_ram[9945] = 8'h00;
    ff_ram[9946] = 8'h00;
    ff_ram[9947] = 8'h00;
    ff_ram[9948] = 8'h00;
    ff_ram[9949] = 8'h00;
    ff_ram[9950] = 8'h00;
    ff_ram[9951] = 8'h00;
    ff_ram[9952] = 8'h00;
    ff_ram[9953] = 8'h00;
    ff_ram[9954] = 8'h00;
    ff_ram[9955] = 8'h00;
    ff_ram[9956] = 8'h00;
    ff_ram[9957] = 8'h00;
    ff_ram[9958] = 8'h00;
    ff_ram[9959] = 8'h00;
    ff_ram[9960] = 8'h00;
    ff_ram[9961] = 8'h00;
    ff_ram[9962] = 8'h00;
    ff_ram[9963] = 8'h00;
    ff_ram[9964] = 8'h00;
    ff_ram[9965] = 8'h00;
    ff_ram[9966] = 8'h00;
    ff_ram[9967] = 8'h00;
    ff_ram[9968] = 8'h00;
    ff_ram[9969] = 8'h00;
    ff_ram[9970] = 8'h00;
    ff_ram[9971] = 8'h00;
    ff_ram[9972] = 8'h00;
    ff_ram[9973] = 8'h00;
    ff_ram[9974] = 8'h00;
    ff_ram[9975] = 8'h00;
    ff_ram[9976] = 8'h00;
    ff_ram[9977] = 8'h00;
    ff_ram[9978] = 8'h00;
    ff_ram[9979] = 8'h00;
    ff_ram[9980] = 8'h00;
    ff_ram[9981] = 8'h00;
    ff_ram[9982] = 8'h00;
    ff_ram[9983] = 8'h00;
    ff_ram[9984] = 8'h00;
    ff_ram[9985] = 8'h00;
    ff_ram[9986] = 8'h00;
    ff_ram[9987] = 8'h00;
    ff_ram[9988] = 8'h00;
    ff_ram[9989] = 8'h00;
    ff_ram[9990] = 8'h00;
    ff_ram[9991] = 8'h00;
    ff_ram[9992] = 8'h00;
    ff_ram[9993] = 8'h00;
    ff_ram[9994] = 8'h00;
    ff_ram[9995] = 8'h00;
    ff_ram[9996] = 8'h00;
    ff_ram[9997] = 8'h00;
    ff_ram[9998] = 8'h00;
    ff_ram[9999] = 8'h00;
    ff_ram[10000] = 8'h00;
    ff_ram[10001] = 8'h00;
    ff_ram[10002] = 8'h00;
    ff_ram[10003] = 8'h00;
    ff_ram[10004] = 8'h00;
    ff_ram[10005] = 8'h00;
    ff_ram[10006] = 8'h00;
    ff_ram[10007] = 8'h00;
    ff_ram[10008] = 8'h00;
    ff_ram[10009] = 8'h00;
    ff_ram[10010] = 8'h00;
    ff_ram[10011] = 8'h00;
    ff_ram[10012] = 8'h00;
    ff_ram[10013] = 8'h00;
    ff_ram[10014] = 8'h00;
    ff_ram[10015] = 8'h00;
    ff_ram[10016] = 8'h00;
    ff_ram[10017] = 8'h00;
    ff_ram[10018] = 8'h00;
    ff_ram[10019] = 8'h00;
    ff_ram[10020] = 8'h00;
    ff_ram[10021] = 8'h00;
    ff_ram[10022] = 8'h00;
    ff_ram[10023] = 8'h00;
    ff_ram[10024] = 8'h00;
    ff_ram[10025] = 8'h00;
    ff_ram[10026] = 8'h00;
    ff_ram[10027] = 8'h00;
    ff_ram[10028] = 8'h00;
    ff_ram[10029] = 8'h00;
    ff_ram[10030] = 8'h00;
    ff_ram[10031] = 8'h00;
    ff_ram[10032] = 8'h00;
    ff_ram[10033] = 8'h00;
    ff_ram[10034] = 8'h00;
    ff_ram[10035] = 8'h00;
    ff_ram[10036] = 8'h00;
    ff_ram[10037] = 8'h00;
    ff_ram[10038] = 8'h00;
    ff_ram[10039] = 8'h00;
    ff_ram[10040] = 8'h00;
    ff_ram[10041] = 8'h00;
    ff_ram[10042] = 8'h00;
    ff_ram[10043] = 8'h00;
    ff_ram[10044] = 8'h00;
    ff_ram[10045] = 8'h00;
    ff_ram[10046] = 8'h00;
    ff_ram[10047] = 8'h00;
    ff_ram[10048] = 8'h00;
    ff_ram[10049] = 8'h00;
    ff_ram[10050] = 8'h00;
    ff_ram[10051] = 8'h00;
    ff_ram[10052] = 8'h00;
    ff_ram[10053] = 8'h00;
    ff_ram[10054] = 8'h00;
    ff_ram[10055] = 8'h00;
    ff_ram[10056] = 8'h00;
    ff_ram[10057] = 8'h00;
    ff_ram[10058] = 8'h00;
    ff_ram[10059] = 8'h00;
    ff_ram[10060] = 8'h00;
    ff_ram[10061] = 8'h00;
    ff_ram[10062] = 8'h00;
    ff_ram[10063] = 8'h00;
    ff_ram[10064] = 8'h00;
    ff_ram[10065] = 8'h00;
    ff_ram[10066] = 8'h00;
    ff_ram[10067] = 8'h00;
    ff_ram[10068] = 8'h00;
    ff_ram[10069] = 8'h00;
    ff_ram[10070] = 8'h00;
    ff_ram[10071] = 8'h00;
    ff_ram[10072] = 8'h00;
    ff_ram[10073] = 8'h00;
    ff_ram[10074] = 8'h00;
    ff_ram[10075] = 8'h00;
    ff_ram[10076] = 8'h00;
    ff_ram[10077] = 8'h00;
    ff_ram[10078] = 8'h00;
    ff_ram[10079] = 8'h00;
    ff_ram[10080] = 8'h00;
    ff_ram[10081] = 8'h00;
    ff_ram[10082] = 8'h00;
    ff_ram[10083] = 8'h00;
    ff_ram[10084] = 8'h00;
    ff_ram[10085] = 8'h00;
    ff_ram[10086] = 8'h00;
    ff_ram[10087] = 8'h00;
    ff_ram[10088] = 8'h00;
    ff_ram[10089] = 8'h00;
    ff_ram[10090] = 8'h00;
    ff_ram[10091] = 8'h00;
    ff_ram[10092] = 8'h00;
    ff_ram[10093] = 8'h00;
    ff_ram[10094] = 8'h00;
    ff_ram[10095] = 8'h00;
    ff_ram[10096] = 8'h00;
    ff_ram[10097] = 8'h00;
    ff_ram[10098] = 8'h00;
    ff_ram[10099] = 8'h00;
    ff_ram[10100] = 8'h00;
    ff_ram[10101] = 8'h00;
    ff_ram[10102] = 8'h00;
    ff_ram[10103] = 8'h00;
    ff_ram[10104] = 8'h00;
    ff_ram[10105] = 8'h00;
    ff_ram[10106] = 8'h00;
    ff_ram[10107] = 8'h00;
    ff_ram[10108] = 8'h00;
    ff_ram[10109] = 8'h00;
    ff_ram[10110] = 8'h00;
    ff_ram[10111] = 8'h00;
    ff_ram[10112] = 8'h00;
    ff_ram[10113] = 8'h00;
    ff_ram[10114] = 8'h00;
    ff_ram[10115] = 8'h00;
    ff_ram[10116] = 8'h00;
    ff_ram[10117] = 8'h00;
    ff_ram[10118] = 8'h00;
    ff_ram[10119] = 8'h00;
    ff_ram[10120] = 8'h00;
    ff_ram[10121] = 8'h00;
    ff_ram[10122] = 8'h00;
    ff_ram[10123] = 8'h00;
    ff_ram[10124] = 8'h00;
    ff_ram[10125] = 8'h00;
    ff_ram[10126] = 8'h00;
    ff_ram[10127] = 8'h00;
    ff_ram[10128] = 8'h00;
    ff_ram[10129] = 8'h00;
    ff_ram[10130] = 8'h00;
    ff_ram[10131] = 8'h00;
    ff_ram[10132] = 8'h00;
    ff_ram[10133] = 8'h00;
    ff_ram[10134] = 8'h00;
    ff_ram[10135] = 8'h00;
    ff_ram[10136] = 8'h00;
    ff_ram[10137] = 8'h00;
    ff_ram[10138] = 8'h00;
    ff_ram[10139] = 8'h00;
    ff_ram[10140] = 8'h00;
    ff_ram[10141] = 8'h00;
    ff_ram[10142] = 8'h00;
    ff_ram[10143] = 8'h00;
    ff_ram[10144] = 8'h00;
    ff_ram[10145] = 8'h00;
    ff_ram[10146] = 8'h00;
    ff_ram[10147] = 8'h00;
    ff_ram[10148] = 8'h00;
    ff_ram[10149] = 8'h00;
    ff_ram[10150] = 8'h00;
    ff_ram[10151] = 8'h00;
    ff_ram[10152] = 8'h00;
    ff_ram[10153] = 8'h00;
    ff_ram[10154] = 8'h00;
    ff_ram[10155] = 8'h00;
    ff_ram[10156] = 8'h00;
    ff_ram[10157] = 8'h00;
    ff_ram[10158] = 8'h00;
    ff_ram[10159] = 8'h00;
    ff_ram[10160] = 8'h00;
    ff_ram[10161] = 8'h00;
    ff_ram[10162] = 8'h00;
    ff_ram[10163] = 8'h00;
    ff_ram[10164] = 8'h00;
    ff_ram[10165] = 8'h00;
    ff_ram[10166] = 8'h00;
    ff_ram[10167] = 8'h00;
    ff_ram[10168] = 8'h00;
    ff_ram[10169] = 8'h00;
    ff_ram[10170] = 8'h00;
    ff_ram[10171] = 8'h00;
    ff_ram[10172] = 8'h00;
    ff_ram[10173] = 8'h00;
    ff_ram[10174] = 8'h00;
    ff_ram[10175] = 8'h00;
    ff_ram[10176] = 8'h00;
    ff_ram[10177] = 8'h00;
    ff_ram[10178] = 8'h00;
    ff_ram[10179] = 8'h00;
    ff_ram[10180] = 8'h00;
    ff_ram[10181] = 8'h00;
    ff_ram[10182] = 8'h00;
    ff_ram[10183] = 8'h00;
    ff_ram[10184] = 8'h00;
    ff_ram[10185] = 8'h00;
    ff_ram[10186] = 8'h00;
    ff_ram[10187] = 8'h00;
    ff_ram[10188] = 8'h00;
    ff_ram[10189] = 8'h00;
    ff_ram[10190] = 8'h00;
    ff_ram[10191] = 8'h00;
    ff_ram[10192] = 8'h00;
    ff_ram[10193] = 8'h00;
    ff_ram[10194] = 8'h00;
    ff_ram[10195] = 8'h00;
    ff_ram[10196] = 8'h00;
    ff_ram[10197] = 8'h00;
    ff_ram[10198] = 8'h00;
    ff_ram[10199] = 8'h00;
    ff_ram[10200] = 8'h00;
    ff_ram[10201] = 8'h00;
    ff_ram[10202] = 8'h00;
    ff_ram[10203] = 8'h00;
    ff_ram[10204] = 8'h00;
    ff_ram[10205] = 8'h00;
    ff_ram[10206] = 8'h00;
    ff_ram[10207] = 8'h00;
    ff_ram[10208] = 8'h00;
    ff_ram[10209] = 8'h00;
    ff_ram[10210] = 8'h00;
    ff_ram[10211] = 8'h00;
    ff_ram[10212] = 8'h00;
    ff_ram[10213] = 8'h00;
    ff_ram[10214] = 8'h00;
    ff_ram[10215] = 8'h00;
    ff_ram[10216] = 8'h00;
    ff_ram[10217] = 8'h00;
    ff_ram[10218] = 8'h00;
    ff_ram[10219] = 8'h00;
    ff_ram[10220] = 8'h00;
    ff_ram[10221] = 8'h00;
    ff_ram[10222] = 8'h00;
    ff_ram[10223] = 8'h00;
    ff_ram[10224] = 8'h00;
    ff_ram[10225] = 8'h00;
    ff_ram[10226] = 8'h00;
    ff_ram[10227] = 8'h00;
    ff_ram[10228] = 8'h00;
    ff_ram[10229] = 8'h00;
    ff_ram[10230] = 8'h00;
    ff_ram[10231] = 8'h00;
    ff_ram[10232] = 8'h00;
    ff_ram[10233] = 8'h00;
    ff_ram[10234] = 8'h00;
    ff_ram[10235] = 8'h00;
    ff_ram[10236] = 8'h00;
    ff_ram[10237] = 8'h00;
    ff_ram[10238] = 8'h00;
    ff_ram[10239] = 8'h00;
    ff_ram[10240] = 8'h00;
    ff_ram[10241] = 8'h00;
    ff_ram[10242] = 8'h00;
    ff_ram[10243] = 8'h00;
    ff_ram[10244] = 8'h00;
    ff_ram[10245] = 8'h00;
    ff_ram[10246] = 8'h00;
    ff_ram[10247] = 8'h00;
    ff_ram[10248] = 8'h00;
    ff_ram[10249] = 8'h00;
    ff_ram[10250] = 8'h00;
    ff_ram[10251] = 8'h00;
    ff_ram[10252] = 8'h00;
    ff_ram[10253] = 8'h00;
    ff_ram[10254] = 8'h00;
    ff_ram[10255] = 8'h00;
    ff_ram[10256] = 8'h00;
    ff_ram[10257] = 8'h00;
    ff_ram[10258] = 8'h00;
    ff_ram[10259] = 8'h00;
    ff_ram[10260] = 8'h00;
    ff_ram[10261] = 8'h00;
    ff_ram[10262] = 8'h00;
    ff_ram[10263] = 8'h00;
    ff_ram[10264] = 8'h00;
    ff_ram[10265] = 8'h00;
    ff_ram[10266] = 8'h00;
    ff_ram[10267] = 8'h00;
    ff_ram[10268] = 8'h00;
    ff_ram[10269] = 8'h00;
    ff_ram[10270] = 8'h00;
    ff_ram[10271] = 8'h00;
    ff_ram[10272] = 8'h00;
    ff_ram[10273] = 8'h00;
    ff_ram[10274] = 8'h00;
    ff_ram[10275] = 8'h00;
    ff_ram[10276] = 8'h00;
    ff_ram[10277] = 8'h00;
    ff_ram[10278] = 8'h00;
    ff_ram[10279] = 8'h00;
    ff_ram[10280] = 8'h00;
    ff_ram[10281] = 8'h00;
    ff_ram[10282] = 8'h00;
    ff_ram[10283] = 8'h00;
    ff_ram[10284] = 8'h00;
    ff_ram[10285] = 8'h00;
    ff_ram[10286] = 8'h00;
    ff_ram[10287] = 8'h00;
    ff_ram[10288] = 8'h00;
    ff_ram[10289] = 8'h00;
    ff_ram[10290] = 8'h00;
    ff_ram[10291] = 8'h00;
    ff_ram[10292] = 8'h00;
    ff_ram[10293] = 8'h00;
    ff_ram[10294] = 8'h00;
    ff_ram[10295] = 8'h00;
    ff_ram[10296] = 8'h00;
    ff_ram[10297] = 8'h00;
    ff_ram[10298] = 8'h00;
    ff_ram[10299] = 8'h00;
    ff_ram[10300] = 8'h00;
    ff_ram[10301] = 8'h00;
    ff_ram[10302] = 8'h00;
    ff_ram[10303] = 8'h00;
    ff_ram[10304] = 8'h00;
    ff_ram[10305] = 8'h00;
    ff_ram[10306] = 8'h00;
    ff_ram[10307] = 8'h00;
    ff_ram[10308] = 8'h00;
    ff_ram[10309] = 8'h00;
    ff_ram[10310] = 8'h00;
    ff_ram[10311] = 8'h00;
    ff_ram[10312] = 8'h00;
    ff_ram[10313] = 8'h00;
    ff_ram[10314] = 8'h00;
    ff_ram[10315] = 8'h00;
    ff_ram[10316] = 8'h00;
    ff_ram[10317] = 8'h00;
    ff_ram[10318] = 8'h00;
    ff_ram[10319] = 8'h00;
    ff_ram[10320] = 8'h00;
    ff_ram[10321] = 8'h00;
    ff_ram[10322] = 8'h00;
    ff_ram[10323] = 8'h00;
    ff_ram[10324] = 8'h00;
    ff_ram[10325] = 8'h00;
    ff_ram[10326] = 8'h00;
    ff_ram[10327] = 8'h00;
    ff_ram[10328] = 8'h00;
    ff_ram[10329] = 8'h00;
    ff_ram[10330] = 8'h00;
    ff_ram[10331] = 8'h00;
    ff_ram[10332] = 8'h00;
    ff_ram[10333] = 8'h00;
    ff_ram[10334] = 8'h00;
    ff_ram[10335] = 8'h00;
    ff_ram[10336] = 8'h00;
    ff_ram[10337] = 8'h00;
    ff_ram[10338] = 8'h00;
    ff_ram[10339] = 8'h00;
    ff_ram[10340] = 8'h00;
    ff_ram[10341] = 8'h00;
    ff_ram[10342] = 8'h00;
    ff_ram[10343] = 8'h00;
    ff_ram[10344] = 8'h00;
    ff_ram[10345] = 8'h00;
    ff_ram[10346] = 8'h00;
    ff_ram[10347] = 8'h00;
    ff_ram[10348] = 8'h00;
    ff_ram[10349] = 8'h00;
    ff_ram[10350] = 8'h00;
    ff_ram[10351] = 8'h00;
    ff_ram[10352] = 8'h00;
    ff_ram[10353] = 8'h00;
    ff_ram[10354] = 8'h00;
    ff_ram[10355] = 8'h00;
    ff_ram[10356] = 8'h00;
    ff_ram[10357] = 8'h00;
    ff_ram[10358] = 8'h00;
    ff_ram[10359] = 8'h00;
    ff_ram[10360] = 8'h00;
    ff_ram[10361] = 8'h00;
    ff_ram[10362] = 8'h00;
    ff_ram[10363] = 8'h00;
    ff_ram[10364] = 8'h00;
    ff_ram[10365] = 8'h00;
    ff_ram[10366] = 8'h00;
    ff_ram[10367] = 8'h00;
    ff_ram[10368] = 8'h00;
    ff_ram[10369] = 8'h00;
    ff_ram[10370] = 8'h00;
    ff_ram[10371] = 8'h00;
    ff_ram[10372] = 8'h00;
    ff_ram[10373] = 8'h00;
    ff_ram[10374] = 8'h00;
    ff_ram[10375] = 8'h00;
    ff_ram[10376] = 8'h00;
    ff_ram[10377] = 8'h00;
    ff_ram[10378] = 8'h00;
    ff_ram[10379] = 8'h00;
    ff_ram[10380] = 8'h00;
    ff_ram[10381] = 8'h00;
    ff_ram[10382] = 8'h00;
    ff_ram[10383] = 8'h00;
    ff_ram[10384] = 8'h00;
    ff_ram[10385] = 8'h00;
    ff_ram[10386] = 8'h00;
    ff_ram[10387] = 8'h00;
    ff_ram[10388] = 8'h00;
    ff_ram[10389] = 8'h00;
    ff_ram[10390] = 8'h00;
    ff_ram[10391] = 8'h00;
    ff_ram[10392] = 8'h00;
    ff_ram[10393] = 8'h00;
    ff_ram[10394] = 8'h00;
    ff_ram[10395] = 8'h00;
    ff_ram[10396] = 8'h00;
    ff_ram[10397] = 8'h00;
    ff_ram[10398] = 8'h00;
    ff_ram[10399] = 8'h00;
    ff_ram[10400] = 8'h00;
    ff_ram[10401] = 8'h00;
    ff_ram[10402] = 8'h00;
    ff_ram[10403] = 8'h00;
    ff_ram[10404] = 8'h00;
    ff_ram[10405] = 8'h00;
    ff_ram[10406] = 8'h00;
    ff_ram[10407] = 8'h00;
    ff_ram[10408] = 8'h00;
    ff_ram[10409] = 8'h00;
    ff_ram[10410] = 8'h00;
    ff_ram[10411] = 8'h00;
    ff_ram[10412] = 8'h00;
    ff_ram[10413] = 8'h00;
    ff_ram[10414] = 8'h00;
    ff_ram[10415] = 8'h00;
    ff_ram[10416] = 8'h00;
    ff_ram[10417] = 8'h00;
    ff_ram[10418] = 8'h00;
    ff_ram[10419] = 8'h00;
    ff_ram[10420] = 8'h00;
    ff_ram[10421] = 8'h00;
    ff_ram[10422] = 8'h00;
    ff_ram[10423] = 8'h00;
    ff_ram[10424] = 8'h00;
    ff_ram[10425] = 8'h00;
    ff_ram[10426] = 8'h00;
    ff_ram[10427] = 8'h00;
    ff_ram[10428] = 8'h00;
    ff_ram[10429] = 8'h00;
    ff_ram[10430] = 8'h00;
    ff_ram[10431] = 8'h00;
    ff_ram[10432] = 8'h00;
    ff_ram[10433] = 8'h00;
    ff_ram[10434] = 8'h00;
    ff_ram[10435] = 8'h00;
    ff_ram[10436] = 8'h00;
    ff_ram[10437] = 8'h00;
    ff_ram[10438] = 8'h00;
    ff_ram[10439] = 8'h00;
    ff_ram[10440] = 8'h00;
    ff_ram[10441] = 8'h00;
    ff_ram[10442] = 8'h00;
    ff_ram[10443] = 8'h00;
    ff_ram[10444] = 8'h00;
    ff_ram[10445] = 8'h00;
    ff_ram[10446] = 8'h00;
    ff_ram[10447] = 8'h00;
    ff_ram[10448] = 8'h00;
    ff_ram[10449] = 8'h00;
    ff_ram[10450] = 8'h00;
    ff_ram[10451] = 8'h00;
    ff_ram[10452] = 8'h00;
    ff_ram[10453] = 8'h00;
    ff_ram[10454] = 8'h00;
    ff_ram[10455] = 8'h00;
    ff_ram[10456] = 8'h00;
    ff_ram[10457] = 8'h00;
    ff_ram[10458] = 8'h00;
    ff_ram[10459] = 8'h00;
    ff_ram[10460] = 8'h00;
    ff_ram[10461] = 8'h00;
    ff_ram[10462] = 8'h00;
    ff_ram[10463] = 8'h00;
    ff_ram[10464] = 8'h00;
    ff_ram[10465] = 8'h00;
    ff_ram[10466] = 8'h00;
    ff_ram[10467] = 8'h00;
    ff_ram[10468] = 8'h00;
    ff_ram[10469] = 8'h00;
    ff_ram[10470] = 8'h00;
    ff_ram[10471] = 8'h00;
    ff_ram[10472] = 8'h00;
    ff_ram[10473] = 8'h00;
    ff_ram[10474] = 8'h00;
    ff_ram[10475] = 8'h00;
    ff_ram[10476] = 8'h00;
    ff_ram[10477] = 8'h00;
    ff_ram[10478] = 8'h00;
    ff_ram[10479] = 8'h00;
    ff_ram[10480] = 8'h00;
    ff_ram[10481] = 8'h00;
    ff_ram[10482] = 8'h00;
    ff_ram[10483] = 8'h00;
    ff_ram[10484] = 8'h00;
    ff_ram[10485] = 8'h00;
    ff_ram[10486] = 8'h00;
    ff_ram[10487] = 8'h00;
    ff_ram[10488] = 8'h00;
    ff_ram[10489] = 8'h00;
    ff_ram[10490] = 8'h00;
    ff_ram[10491] = 8'h00;
    ff_ram[10492] = 8'h00;
    ff_ram[10493] = 8'h00;
    ff_ram[10494] = 8'h00;
    ff_ram[10495] = 8'h00;
    ff_ram[10496] = 8'h00;
    ff_ram[10497] = 8'h00;
    ff_ram[10498] = 8'h00;
    ff_ram[10499] = 8'h00;
    ff_ram[10500] = 8'h00;
    ff_ram[10501] = 8'h00;
    ff_ram[10502] = 8'h00;
    ff_ram[10503] = 8'h00;
    ff_ram[10504] = 8'h00;
    ff_ram[10505] = 8'h00;
    ff_ram[10506] = 8'h00;
    ff_ram[10507] = 8'h00;
    ff_ram[10508] = 8'h00;
    ff_ram[10509] = 8'h00;
    ff_ram[10510] = 8'h00;
    ff_ram[10511] = 8'h00;
    ff_ram[10512] = 8'h00;
    ff_ram[10513] = 8'h00;
    ff_ram[10514] = 8'h00;
    ff_ram[10515] = 8'h00;
    ff_ram[10516] = 8'h00;
    ff_ram[10517] = 8'h00;
    ff_ram[10518] = 8'h00;
    ff_ram[10519] = 8'h00;
    ff_ram[10520] = 8'h00;
    ff_ram[10521] = 8'h00;
    ff_ram[10522] = 8'h00;
    ff_ram[10523] = 8'h00;
    ff_ram[10524] = 8'h00;
    ff_ram[10525] = 8'h00;
    ff_ram[10526] = 8'h00;
    ff_ram[10527] = 8'h00;
    ff_ram[10528] = 8'h00;
    ff_ram[10529] = 8'h00;
    ff_ram[10530] = 8'h00;
    ff_ram[10531] = 8'h00;
    ff_ram[10532] = 8'h00;
    ff_ram[10533] = 8'h00;
    ff_ram[10534] = 8'h00;
    ff_ram[10535] = 8'h00;
    ff_ram[10536] = 8'h00;
    ff_ram[10537] = 8'h00;
    ff_ram[10538] = 8'h00;
    ff_ram[10539] = 8'h00;
    ff_ram[10540] = 8'h00;
    ff_ram[10541] = 8'h00;
    ff_ram[10542] = 8'h00;
    ff_ram[10543] = 8'h00;
    ff_ram[10544] = 8'h00;
    ff_ram[10545] = 8'h00;
    ff_ram[10546] = 8'h00;
    ff_ram[10547] = 8'h00;
    ff_ram[10548] = 8'h00;
    ff_ram[10549] = 8'h00;
    ff_ram[10550] = 8'h00;
    ff_ram[10551] = 8'h00;
    ff_ram[10552] = 8'h00;
    ff_ram[10553] = 8'h00;
    ff_ram[10554] = 8'h00;
    ff_ram[10555] = 8'h00;
    ff_ram[10556] = 8'h00;
    ff_ram[10557] = 8'h00;
    ff_ram[10558] = 8'h00;
    ff_ram[10559] = 8'h00;
    ff_ram[10560] = 8'h00;
    ff_ram[10561] = 8'h00;
    ff_ram[10562] = 8'h00;
    ff_ram[10563] = 8'h00;
    ff_ram[10564] = 8'h00;
    ff_ram[10565] = 8'h00;
    ff_ram[10566] = 8'h00;
    ff_ram[10567] = 8'h00;
    ff_ram[10568] = 8'h00;
    ff_ram[10569] = 8'h00;
    ff_ram[10570] = 8'h00;
    ff_ram[10571] = 8'h00;
    ff_ram[10572] = 8'h00;
    ff_ram[10573] = 8'h00;
    ff_ram[10574] = 8'h00;
    ff_ram[10575] = 8'h00;
    ff_ram[10576] = 8'h00;
    ff_ram[10577] = 8'h00;
    ff_ram[10578] = 8'h00;
    ff_ram[10579] = 8'h00;
    ff_ram[10580] = 8'h00;
    ff_ram[10581] = 8'h00;
    ff_ram[10582] = 8'h00;
    ff_ram[10583] = 8'h00;
    ff_ram[10584] = 8'h00;
    ff_ram[10585] = 8'h00;
    ff_ram[10586] = 8'h00;
    ff_ram[10587] = 8'h00;
    ff_ram[10588] = 8'h00;
    ff_ram[10589] = 8'h00;
    ff_ram[10590] = 8'h00;
    ff_ram[10591] = 8'h00;
    ff_ram[10592] = 8'h00;
    ff_ram[10593] = 8'h00;
    ff_ram[10594] = 8'h00;
    ff_ram[10595] = 8'h00;
    ff_ram[10596] = 8'h00;
    ff_ram[10597] = 8'h00;
    ff_ram[10598] = 8'h00;
    ff_ram[10599] = 8'h00;
    ff_ram[10600] = 8'h00;
    ff_ram[10601] = 8'h00;
    ff_ram[10602] = 8'h00;
    ff_ram[10603] = 8'h00;
    ff_ram[10604] = 8'h00;
    ff_ram[10605] = 8'h00;
    ff_ram[10606] = 8'h00;
    ff_ram[10607] = 8'h00;
    ff_ram[10608] = 8'h00;
    ff_ram[10609] = 8'h00;
    ff_ram[10610] = 8'h00;
    ff_ram[10611] = 8'h00;
    ff_ram[10612] = 8'h00;
    ff_ram[10613] = 8'h00;
    ff_ram[10614] = 8'h00;
    ff_ram[10615] = 8'h00;
    ff_ram[10616] = 8'h00;
    ff_ram[10617] = 8'h00;
    ff_ram[10618] = 8'h00;
    ff_ram[10619] = 8'h00;
    ff_ram[10620] = 8'h00;
    ff_ram[10621] = 8'h00;
    ff_ram[10622] = 8'h00;
    ff_ram[10623] = 8'h00;
    ff_ram[10624] = 8'h00;
    ff_ram[10625] = 8'h00;
    ff_ram[10626] = 8'h00;
    ff_ram[10627] = 8'h00;
    ff_ram[10628] = 8'h00;
    ff_ram[10629] = 8'h00;
    ff_ram[10630] = 8'h00;
    ff_ram[10631] = 8'h00;
    ff_ram[10632] = 8'h00;
    ff_ram[10633] = 8'h00;
    ff_ram[10634] = 8'h00;
    ff_ram[10635] = 8'h00;
    ff_ram[10636] = 8'h00;
    ff_ram[10637] = 8'h00;
    ff_ram[10638] = 8'h00;
    ff_ram[10639] = 8'h00;
    ff_ram[10640] = 8'h00;
    ff_ram[10641] = 8'h00;
    ff_ram[10642] = 8'h00;
    ff_ram[10643] = 8'h00;
    ff_ram[10644] = 8'h00;
    ff_ram[10645] = 8'h00;
    ff_ram[10646] = 8'h00;
    ff_ram[10647] = 8'h00;
    ff_ram[10648] = 8'h00;
    ff_ram[10649] = 8'h00;
    ff_ram[10650] = 8'h00;
    ff_ram[10651] = 8'h00;
    ff_ram[10652] = 8'h00;
    ff_ram[10653] = 8'h00;
    ff_ram[10654] = 8'h00;
    ff_ram[10655] = 8'h00;
    ff_ram[10656] = 8'h00;
    ff_ram[10657] = 8'h00;
    ff_ram[10658] = 8'h00;
    ff_ram[10659] = 8'h00;
    ff_ram[10660] = 8'h00;
    ff_ram[10661] = 8'h00;
    ff_ram[10662] = 8'h00;
    ff_ram[10663] = 8'h00;
    ff_ram[10664] = 8'h00;
    ff_ram[10665] = 8'h00;
    ff_ram[10666] = 8'h00;
    ff_ram[10667] = 8'h00;
    ff_ram[10668] = 8'h00;
    ff_ram[10669] = 8'h00;
    ff_ram[10670] = 8'h00;
    ff_ram[10671] = 8'h00;
    ff_ram[10672] = 8'h00;
    ff_ram[10673] = 8'h00;
    ff_ram[10674] = 8'h00;
    ff_ram[10675] = 8'h00;
    ff_ram[10676] = 8'h00;
    ff_ram[10677] = 8'h00;
    ff_ram[10678] = 8'h00;
    ff_ram[10679] = 8'h00;
    ff_ram[10680] = 8'h00;
    ff_ram[10681] = 8'h00;
    ff_ram[10682] = 8'h00;
    ff_ram[10683] = 8'h00;
    ff_ram[10684] = 8'h00;
    ff_ram[10685] = 8'h00;
    ff_ram[10686] = 8'h00;
    ff_ram[10687] = 8'h00;
    ff_ram[10688] = 8'h00;
    ff_ram[10689] = 8'h00;
    ff_ram[10690] = 8'h00;
    ff_ram[10691] = 8'h00;
    ff_ram[10692] = 8'h00;
    ff_ram[10693] = 8'h00;
    ff_ram[10694] = 8'h00;
    ff_ram[10695] = 8'h00;
    ff_ram[10696] = 8'h00;
    ff_ram[10697] = 8'h00;
    ff_ram[10698] = 8'h00;
    ff_ram[10699] = 8'h00;
    ff_ram[10700] = 8'h00;
    ff_ram[10701] = 8'h00;
    ff_ram[10702] = 8'h00;
    ff_ram[10703] = 8'h00;
    ff_ram[10704] = 8'h00;
    ff_ram[10705] = 8'h00;
    ff_ram[10706] = 8'h00;
    ff_ram[10707] = 8'h00;
    ff_ram[10708] = 8'h00;
    ff_ram[10709] = 8'h00;
    ff_ram[10710] = 8'h00;
    ff_ram[10711] = 8'h00;
    ff_ram[10712] = 8'h00;
    ff_ram[10713] = 8'h00;
    ff_ram[10714] = 8'h00;
    ff_ram[10715] = 8'h00;
    ff_ram[10716] = 8'h00;
    ff_ram[10717] = 8'h00;
    ff_ram[10718] = 8'h00;
    ff_ram[10719] = 8'h00;
    ff_ram[10720] = 8'h00;
    ff_ram[10721] = 8'h00;
    ff_ram[10722] = 8'h00;
    ff_ram[10723] = 8'h00;
    ff_ram[10724] = 8'h00;
    ff_ram[10725] = 8'h00;
    ff_ram[10726] = 8'h00;
    ff_ram[10727] = 8'h00;
    ff_ram[10728] = 8'h00;
    ff_ram[10729] = 8'h00;
    ff_ram[10730] = 8'h00;
    ff_ram[10731] = 8'h00;
    ff_ram[10732] = 8'h00;
    ff_ram[10733] = 8'h00;
    ff_ram[10734] = 8'h00;
    ff_ram[10735] = 8'h00;
    ff_ram[10736] = 8'h00;
    ff_ram[10737] = 8'h00;
    ff_ram[10738] = 8'h00;
    ff_ram[10739] = 8'h00;
    ff_ram[10740] = 8'h00;
    ff_ram[10741] = 8'h00;
    ff_ram[10742] = 8'h00;
    ff_ram[10743] = 8'h00;
    ff_ram[10744] = 8'h00;
    ff_ram[10745] = 8'h00;
    ff_ram[10746] = 8'h00;
    ff_ram[10747] = 8'h00;
    ff_ram[10748] = 8'h00;
    ff_ram[10749] = 8'h00;
    ff_ram[10750] = 8'h00;
    ff_ram[10751] = 8'h00;
    ff_ram[10752] = 8'h00;
    ff_ram[10753] = 8'h00;
    ff_ram[10754] = 8'h00;
    ff_ram[10755] = 8'h00;
    ff_ram[10756] = 8'h00;
    ff_ram[10757] = 8'h00;
    ff_ram[10758] = 8'h00;
    ff_ram[10759] = 8'h00;
    ff_ram[10760] = 8'h00;
    ff_ram[10761] = 8'h00;
    ff_ram[10762] = 8'h00;
    ff_ram[10763] = 8'h00;
    ff_ram[10764] = 8'h00;
    ff_ram[10765] = 8'h00;
    ff_ram[10766] = 8'h00;
    ff_ram[10767] = 8'h00;
    ff_ram[10768] = 8'h00;
    ff_ram[10769] = 8'h00;
    ff_ram[10770] = 8'h00;
    ff_ram[10771] = 8'h00;
    ff_ram[10772] = 8'h00;
    ff_ram[10773] = 8'h00;
    ff_ram[10774] = 8'h00;
    ff_ram[10775] = 8'h00;
    ff_ram[10776] = 8'h00;
    ff_ram[10777] = 8'h00;
    ff_ram[10778] = 8'h00;
    ff_ram[10779] = 8'h00;
    ff_ram[10780] = 8'h00;
    ff_ram[10781] = 8'h00;
    ff_ram[10782] = 8'h00;
    ff_ram[10783] = 8'h00;
    ff_ram[10784] = 8'h00;
    ff_ram[10785] = 8'h00;
    ff_ram[10786] = 8'h00;
    ff_ram[10787] = 8'h00;
    ff_ram[10788] = 8'h00;
    ff_ram[10789] = 8'h00;
    ff_ram[10790] = 8'h00;
    ff_ram[10791] = 8'h00;
    ff_ram[10792] = 8'h00;
    ff_ram[10793] = 8'h00;
    ff_ram[10794] = 8'h00;
    ff_ram[10795] = 8'h00;
    ff_ram[10796] = 8'h00;
    ff_ram[10797] = 8'h00;
    ff_ram[10798] = 8'h00;
    ff_ram[10799] = 8'h00;
    ff_ram[10800] = 8'h00;
    ff_ram[10801] = 8'h00;
    ff_ram[10802] = 8'h00;
    ff_ram[10803] = 8'h00;
    ff_ram[10804] = 8'h00;
    ff_ram[10805] = 8'h00;
    ff_ram[10806] = 8'h00;
    ff_ram[10807] = 8'h00;
    ff_ram[10808] = 8'h00;
    ff_ram[10809] = 8'h00;
    ff_ram[10810] = 8'h00;
    ff_ram[10811] = 8'h00;
    ff_ram[10812] = 8'h00;
    ff_ram[10813] = 8'h00;
    ff_ram[10814] = 8'h00;
    ff_ram[10815] = 8'h00;
    ff_ram[10816] = 8'h00;
    ff_ram[10817] = 8'h00;
    ff_ram[10818] = 8'h00;
    ff_ram[10819] = 8'h00;
    ff_ram[10820] = 8'h00;
    ff_ram[10821] = 8'h00;
    ff_ram[10822] = 8'h00;
    ff_ram[10823] = 8'h00;
    ff_ram[10824] = 8'h00;
    ff_ram[10825] = 8'h00;
    ff_ram[10826] = 8'h00;
    ff_ram[10827] = 8'h00;
    ff_ram[10828] = 8'h00;
    ff_ram[10829] = 8'h00;
    ff_ram[10830] = 8'h00;
    ff_ram[10831] = 8'h00;
    ff_ram[10832] = 8'h00;
    ff_ram[10833] = 8'h00;
    ff_ram[10834] = 8'h00;
    ff_ram[10835] = 8'h00;
    ff_ram[10836] = 8'h00;
    ff_ram[10837] = 8'h00;
    ff_ram[10838] = 8'h00;
    ff_ram[10839] = 8'h00;
    ff_ram[10840] = 8'h00;
    ff_ram[10841] = 8'h00;
    ff_ram[10842] = 8'h00;
    ff_ram[10843] = 8'h00;
    ff_ram[10844] = 8'h00;
    ff_ram[10845] = 8'h00;
    ff_ram[10846] = 8'h00;
    ff_ram[10847] = 8'h00;
    ff_ram[10848] = 8'h00;
    ff_ram[10849] = 8'h00;
    ff_ram[10850] = 8'h00;
    ff_ram[10851] = 8'h00;
    ff_ram[10852] = 8'h00;
    ff_ram[10853] = 8'h00;
    ff_ram[10854] = 8'h00;
    ff_ram[10855] = 8'h00;
    ff_ram[10856] = 8'h00;
    ff_ram[10857] = 8'h00;
    ff_ram[10858] = 8'h00;
    ff_ram[10859] = 8'h00;
    ff_ram[10860] = 8'h00;
    ff_ram[10861] = 8'h00;
    ff_ram[10862] = 8'h00;
    ff_ram[10863] = 8'h00;
    ff_ram[10864] = 8'h00;
    ff_ram[10865] = 8'h00;
    ff_ram[10866] = 8'h00;
    ff_ram[10867] = 8'h00;
    ff_ram[10868] = 8'h00;
    ff_ram[10869] = 8'h00;
    ff_ram[10870] = 8'h00;
    ff_ram[10871] = 8'h00;
    ff_ram[10872] = 8'h00;
    ff_ram[10873] = 8'h00;
    ff_ram[10874] = 8'h00;
    ff_ram[10875] = 8'h00;
    ff_ram[10876] = 8'h00;
    ff_ram[10877] = 8'h00;
    ff_ram[10878] = 8'h00;
    ff_ram[10879] = 8'h00;
    ff_ram[10880] = 8'h00;
    ff_ram[10881] = 8'h00;
    ff_ram[10882] = 8'h00;
    ff_ram[10883] = 8'h00;
    ff_ram[10884] = 8'h00;
    ff_ram[10885] = 8'h00;
    ff_ram[10886] = 8'h00;
    ff_ram[10887] = 8'h00;
    ff_ram[10888] = 8'h00;
    ff_ram[10889] = 8'h00;
    ff_ram[10890] = 8'h00;
    ff_ram[10891] = 8'h00;
    ff_ram[10892] = 8'h00;
    ff_ram[10893] = 8'h00;
    ff_ram[10894] = 8'h00;
    ff_ram[10895] = 8'h00;
    ff_ram[10896] = 8'h00;
    ff_ram[10897] = 8'h00;
    ff_ram[10898] = 8'h00;
    ff_ram[10899] = 8'h00;
    ff_ram[10900] = 8'h00;
    ff_ram[10901] = 8'h00;
    ff_ram[10902] = 8'h00;
    ff_ram[10903] = 8'h00;
    ff_ram[10904] = 8'h00;
    ff_ram[10905] = 8'h00;
    ff_ram[10906] = 8'h00;
    ff_ram[10907] = 8'h00;
    ff_ram[10908] = 8'h00;
    ff_ram[10909] = 8'h00;
    ff_ram[10910] = 8'h00;
    ff_ram[10911] = 8'h00;
    ff_ram[10912] = 8'h00;
    ff_ram[10913] = 8'h00;
    ff_ram[10914] = 8'h00;
    ff_ram[10915] = 8'h00;
    ff_ram[10916] = 8'h00;
    ff_ram[10917] = 8'h00;
    ff_ram[10918] = 8'h00;
    ff_ram[10919] = 8'h00;
    ff_ram[10920] = 8'h00;
    ff_ram[10921] = 8'h00;
    ff_ram[10922] = 8'h00;
    ff_ram[10923] = 8'h00;
    ff_ram[10924] = 8'h00;
    ff_ram[10925] = 8'h00;
    ff_ram[10926] = 8'h00;
    ff_ram[10927] = 8'h00;
    ff_ram[10928] = 8'h00;
    ff_ram[10929] = 8'h00;
    ff_ram[10930] = 8'h00;
    ff_ram[10931] = 8'h00;
    ff_ram[10932] = 8'h00;
    ff_ram[10933] = 8'h00;
    ff_ram[10934] = 8'h00;
    ff_ram[10935] = 8'h00;
    ff_ram[10936] = 8'h00;
    ff_ram[10937] = 8'h00;
    ff_ram[10938] = 8'h00;
    ff_ram[10939] = 8'h00;
    ff_ram[10940] = 8'h00;
    ff_ram[10941] = 8'h00;
    ff_ram[10942] = 8'h00;
    ff_ram[10943] = 8'h00;
    ff_ram[10944] = 8'h00;
    ff_ram[10945] = 8'h00;
    ff_ram[10946] = 8'h00;
    ff_ram[10947] = 8'h00;
    ff_ram[10948] = 8'h00;
    ff_ram[10949] = 8'h00;
    ff_ram[10950] = 8'h00;
    ff_ram[10951] = 8'h00;
    ff_ram[10952] = 8'h00;
    ff_ram[10953] = 8'h00;
    ff_ram[10954] = 8'h00;
    ff_ram[10955] = 8'h00;
    ff_ram[10956] = 8'h00;
    ff_ram[10957] = 8'h00;
    ff_ram[10958] = 8'h00;
    ff_ram[10959] = 8'h00;
    ff_ram[10960] = 8'h00;
    ff_ram[10961] = 8'h00;
    ff_ram[10962] = 8'h00;
    ff_ram[10963] = 8'h00;
    ff_ram[10964] = 8'h00;
    ff_ram[10965] = 8'h00;
    ff_ram[10966] = 8'h00;
    ff_ram[10967] = 8'h00;
    ff_ram[10968] = 8'h00;
    ff_ram[10969] = 8'h00;
    ff_ram[10970] = 8'h00;
    ff_ram[10971] = 8'h00;
    ff_ram[10972] = 8'h00;
    ff_ram[10973] = 8'h00;
    ff_ram[10974] = 8'h00;
    ff_ram[10975] = 8'h00;
    ff_ram[10976] = 8'h00;
    ff_ram[10977] = 8'h00;
    ff_ram[10978] = 8'h00;
    ff_ram[10979] = 8'h00;
    ff_ram[10980] = 8'h00;
    ff_ram[10981] = 8'h00;
    ff_ram[10982] = 8'h00;
    ff_ram[10983] = 8'h00;
    ff_ram[10984] = 8'h00;
    ff_ram[10985] = 8'h00;
    ff_ram[10986] = 8'h00;
    ff_ram[10987] = 8'h00;
    ff_ram[10988] = 8'h00;
    ff_ram[10989] = 8'h00;
    ff_ram[10990] = 8'h00;
    ff_ram[10991] = 8'h00;
    ff_ram[10992] = 8'h00;
    ff_ram[10993] = 8'h00;
    ff_ram[10994] = 8'h00;
    ff_ram[10995] = 8'h00;
    ff_ram[10996] = 8'h00;
    ff_ram[10997] = 8'h00;
    ff_ram[10998] = 8'h00;
    ff_ram[10999] = 8'h00;
    ff_ram[11000] = 8'h00;
    ff_ram[11001] = 8'h00;
    ff_ram[11002] = 8'h00;
    ff_ram[11003] = 8'h00;
    ff_ram[11004] = 8'h00;
    ff_ram[11005] = 8'h00;
    ff_ram[11006] = 8'h00;
    ff_ram[11007] = 8'h00;
    ff_ram[11008] = 8'h00;
    ff_ram[11009] = 8'h00;
    ff_ram[11010] = 8'h00;
    ff_ram[11011] = 8'h00;
    ff_ram[11012] = 8'h00;
    ff_ram[11013] = 8'h00;
    ff_ram[11014] = 8'h00;
    ff_ram[11015] = 8'h00;
    ff_ram[11016] = 8'h00;
    ff_ram[11017] = 8'h00;
    ff_ram[11018] = 8'h00;
    ff_ram[11019] = 8'h00;
    ff_ram[11020] = 8'h00;
    ff_ram[11021] = 8'h00;
    ff_ram[11022] = 8'h00;
    ff_ram[11023] = 8'h00;
    ff_ram[11024] = 8'h00;
    ff_ram[11025] = 8'h00;
    ff_ram[11026] = 8'h00;
    ff_ram[11027] = 8'h00;
    ff_ram[11028] = 8'h00;
    ff_ram[11029] = 8'h00;
    ff_ram[11030] = 8'h00;
    ff_ram[11031] = 8'h00;
    ff_ram[11032] = 8'h00;
    ff_ram[11033] = 8'h00;
    ff_ram[11034] = 8'h00;
    ff_ram[11035] = 8'h00;
    ff_ram[11036] = 8'h00;
    ff_ram[11037] = 8'h00;
    ff_ram[11038] = 8'h00;
    ff_ram[11039] = 8'h00;
    ff_ram[11040] = 8'h00;
    ff_ram[11041] = 8'h00;
    ff_ram[11042] = 8'h00;
    ff_ram[11043] = 8'h00;
    ff_ram[11044] = 8'h00;
    ff_ram[11045] = 8'h00;
    ff_ram[11046] = 8'h00;
    ff_ram[11047] = 8'h00;
    ff_ram[11048] = 8'h00;
    ff_ram[11049] = 8'h00;
    ff_ram[11050] = 8'h00;
    ff_ram[11051] = 8'h00;
    ff_ram[11052] = 8'h00;
    ff_ram[11053] = 8'h00;
    ff_ram[11054] = 8'h00;
    ff_ram[11055] = 8'h00;
    ff_ram[11056] = 8'h00;
    ff_ram[11057] = 8'h00;
    ff_ram[11058] = 8'h00;
    ff_ram[11059] = 8'h00;
    ff_ram[11060] = 8'h00;
    ff_ram[11061] = 8'h00;
    ff_ram[11062] = 8'h00;
    ff_ram[11063] = 8'h00;
    ff_ram[11064] = 8'h00;
    ff_ram[11065] = 8'h00;
    ff_ram[11066] = 8'h00;
    ff_ram[11067] = 8'h00;
    ff_ram[11068] = 8'h00;
    ff_ram[11069] = 8'h00;
    ff_ram[11070] = 8'h00;
    ff_ram[11071] = 8'h00;
    ff_ram[11072] = 8'h00;
    ff_ram[11073] = 8'h00;
    ff_ram[11074] = 8'h00;
    ff_ram[11075] = 8'h00;
    ff_ram[11076] = 8'h00;
    ff_ram[11077] = 8'h00;
    ff_ram[11078] = 8'h00;
    ff_ram[11079] = 8'h00;
    ff_ram[11080] = 8'h00;
    ff_ram[11081] = 8'h00;
    ff_ram[11082] = 8'h00;
    ff_ram[11083] = 8'h00;
    ff_ram[11084] = 8'h00;
    ff_ram[11085] = 8'h00;
    ff_ram[11086] = 8'h00;
    ff_ram[11087] = 8'h00;
    ff_ram[11088] = 8'h00;
    ff_ram[11089] = 8'h00;
    ff_ram[11090] = 8'h00;
    ff_ram[11091] = 8'h00;
    ff_ram[11092] = 8'h00;
    ff_ram[11093] = 8'h00;
    ff_ram[11094] = 8'h00;
    ff_ram[11095] = 8'h00;
    ff_ram[11096] = 8'h00;
    ff_ram[11097] = 8'h00;
    ff_ram[11098] = 8'h00;
    ff_ram[11099] = 8'h00;
    ff_ram[11100] = 8'h00;
    ff_ram[11101] = 8'h00;
    ff_ram[11102] = 8'h00;
    ff_ram[11103] = 8'h00;
    ff_ram[11104] = 8'h00;
    ff_ram[11105] = 8'h00;
    ff_ram[11106] = 8'h00;
    ff_ram[11107] = 8'h00;
    ff_ram[11108] = 8'h00;
    ff_ram[11109] = 8'h00;
    ff_ram[11110] = 8'h00;
    ff_ram[11111] = 8'h00;
    ff_ram[11112] = 8'h00;
    ff_ram[11113] = 8'h00;
    ff_ram[11114] = 8'h00;
    ff_ram[11115] = 8'h00;
    ff_ram[11116] = 8'h00;
    ff_ram[11117] = 8'h00;
    ff_ram[11118] = 8'h00;
    ff_ram[11119] = 8'h00;
    ff_ram[11120] = 8'h00;
    ff_ram[11121] = 8'h00;
    ff_ram[11122] = 8'h00;
    ff_ram[11123] = 8'h00;
    ff_ram[11124] = 8'h00;
    ff_ram[11125] = 8'h00;
    ff_ram[11126] = 8'h00;
    ff_ram[11127] = 8'h00;
    ff_ram[11128] = 8'h00;
    ff_ram[11129] = 8'h00;
    ff_ram[11130] = 8'h00;
    ff_ram[11131] = 8'h00;
    ff_ram[11132] = 8'h00;
    ff_ram[11133] = 8'h00;
    ff_ram[11134] = 8'h00;
    ff_ram[11135] = 8'h00;
    ff_ram[11136] = 8'h00;
    ff_ram[11137] = 8'h00;
    ff_ram[11138] = 8'h00;
    ff_ram[11139] = 8'h00;
    ff_ram[11140] = 8'h00;
    ff_ram[11141] = 8'h00;
    ff_ram[11142] = 8'h00;
    ff_ram[11143] = 8'h00;
    ff_ram[11144] = 8'h00;
    ff_ram[11145] = 8'h00;
    ff_ram[11146] = 8'h00;
    ff_ram[11147] = 8'h00;
    ff_ram[11148] = 8'h00;
    ff_ram[11149] = 8'h00;
    ff_ram[11150] = 8'h00;
    ff_ram[11151] = 8'h00;
    ff_ram[11152] = 8'h00;
    ff_ram[11153] = 8'h00;
    ff_ram[11154] = 8'h00;
    ff_ram[11155] = 8'h00;
    ff_ram[11156] = 8'h00;
    ff_ram[11157] = 8'h00;
    ff_ram[11158] = 8'h00;
    ff_ram[11159] = 8'h00;
    ff_ram[11160] = 8'h00;
    ff_ram[11161] = 8'h00;
    ff_ram[11162] = 8'h00;
    ff_ram[11163] = 8'h00;
    ff_ram[11164] = 8'h00;
    ff_ram[11165] = 8'h00;
    ff_ram[11166] = 8'h00;
    ff_ram[11167] = 8'h00;
    ff_ram[11168] = 8'h00;
    ff_ram[11169] = 8'h00;
    ff_ram[11170] = 8'h00;
    ff_ram[11171] = 8'h00;
    ff_ram[11172] = 8'h00;
    ff_ram[11173] = 8'h00;
    ff_ram[11174] = 8'h00;
    ff_ram[11175] = 8'h00;
    ff_ram[11176] = 8'h00;
    ff_ram[11177] = 8'h00;
    ff_ram[11178] = 8'h00;
    ff_ram[11179] = 8'h00;
    ff_ram[11180] = 8'h00;
    ff_ram[11181] = 8'h00;
    ff_ram[11182] = 8'h00;
    ff_ram[11183] = 8'h00;
    ff_ram[11184] = 8'h00;
    ff_ram[11185] = 8'h00;
    ff_ram[11186] = 8'h00;
    ff_ram[11187] = 8'h00;
    ff_ram[11188] = 8'h00;
    ff_ram[11189] = 8'h00;
    ff_ram[11190] = 8'h00;
    ff_ram[11191] = 8'h00;
    ff_ram[11192] = 8'h00;
    ff_ram[11193] = 8'h00;
    ff_ram[11194] = 8'h00;
    ff_ram[11195] = 8'h00;
    ff_ram[11196] = 8'h00;
    ff_ram[11197] = 8'h00;
    ff_ram[11198] = 8'h00;
    ff_ram[11199] = 8'h00;
    ff_ram[11200] = 8'h00;
    ff_ram[11201] = 8'h00;
    ff_ram[11202] = 8'h00;
    ff_ram[11203] = 8'h00;
    ff_ram[11204] = 8'h00;
    ff_ram[11205] = 8'h00;
    ff_ram[11206] = 8'h00;
    ff_ram[11207] = 8'h00;
    ff_ram[11208] = 8'h00;
    ff_ram[11209] = 8'h00;
    ff_ram[11210] = 8'h00;
    ff_ram[11211] = 8'h00;
    ff_ram[11212] = 8'h00;
    ff_ram[11213] = 8'h00;
    ff_ram[11214] = 8'h00;
    ff_ram[11215] = 8'h00;
    ff_ram[11216] = 8'h00;
    ff_ram[11217] = 8'h00;
    ff_ram[11218] = 8'h00;
    ff_ram[11219] = 8'h00;
    ff_ram[11220] = 8'h00;
    ff_ram[11221] = 8'h00;
    ff_ram[11222] = 8'h00;
    ff_ram[11223] = 8'h00;
    ff_ram[11224] = 8'h00;
    ff_ram[11225] = 8'h00;
    ff_ram[11226] = 8'h00;
    ff_ram[11227] = 8'h00;
    ff_ram[11228] = 8'h00;
    ff_ram[11229] = 8'h00;
    ff_ram[11230] = 8'h00;
    ff_ram[11231] = 8'h00;
    ff_ram[11232] = 8'h00;
    ff_ram[11233] = 8'h00;
    ff_ram[11234] = 8'h00;
    ff_ram[11235] = 8'h00;
    ff_ram[11236] = 8'h00;
    ff_ram[11237] = 8'h00;
    ff_ram[11238] = 8'h00;
    ff_ram[11239] = 8'h00;
    ff_ram[11240] = 8'h00;
    ff_ram[11241] = 8'h00;
    ff_ram[11242] = 8'h00;
    ff_ram[11243] = 8'h00;
    ff_ram[11244] = 8'h00;
    ff_ram[11245] = 8'h00;
    ff_ram[11246] = 8'h00;
    ff_ram[11247] = 8'h00;
    ff_ram[11248] = 8'h00;
    ff_ram[11249] = 8'h00;
    ff_ram[11250] = 8'h00;
    ff_ram[11251] = 8'h00;
    ff_ram[11252] = 8'h00;
    ff_ram[11253] = 8'h00;
    ff_ram[11254] = 8'h00;
    ff_ram[11255] = 8'h00;
    ff_ram[11256] = 8'h00;
    ff_ram[11257] = 8'h00;
    ff_ram[11258] = 8'h00;
    ff_ram[11259] = 8'h00;
    ff_ram[11260] = 8'h00;
    ff_ram[11261] = 8'h00;
    ff_ram[11262] = 8'h00;
    ff_ram[11263] = 8'h00;
    ff_ram[11264] = 8'h00;
    ff_ram[11265] = 8'h00;
    ff_ram[11266] = 8'h00;
    ff_ram[11267] = 8'h00;
    ff_ram[11268] = 8'h00;
    ff_ram[11269] = 8'h00;
    ff_ram[11270] = 8'h00;
    ff_ram[11271] = 8'h00;
    ff_ram[11272] = 8'h00;
    ff_ram[11273] = 8'h00;
    ff_ram[11274] = 8'h00;
    ff_ram[11275] = 8'h00;
    ff_ram[11276] = 8'h00;
    ff_ram[11277] = 8'h00;
    ff_ram[11278] = 8'h00;
    ff_ram[11279] = 8'h00;
    ff_ram[11280] = 8'h00;
    ff_ram[11281] = 8'h00;
    ff_ram[11282] = 8'h00;
    ff_ram[11283] = 8'h00;
    ff_ram[11284] = 8'h00;
    ff_ram[11285] = 8'h00;
    ff_ram[11286] = 8'h00;
    ff_ram[11287] = 8'h00;
    ff_ram[11288] = 8'h00;
    ff_ram[11289] = 8'h00;
    ff_ram[11290] = 8'h00;
    ff_ram[11291] = 8'h00;
    ff_ram[11292] = 8'h00;
    ff_ram[11293] = 8'h00;
    ff_ram[11294] = 8'h00;
    ff_ram[11295] = 8'h00;
    ff_ram[11296] = 8'h00;
    ff_ram[11297] = 8'h00;
    ff_ram[11298] = 8'h00;
    ff_ram[11299] = 8'h00;
    ff_ram[11300] = 8'h00;
    ff_ram[11301] = 8'h00;
    ff_ram[11302] = 8'h00;
    ff_ram[11303] = 8'h00;
    ff_ram[11304] = 8'h00;
    ff_ram[11305] = 8'h00;
    ff_ram[11306] = 8'h00;
    ff_ram[11307] = 8'h00;
    ff_ram[11308] = 8'h00;
    ff_ram[11309] = 8'h00;
    ff_ram[11310] = 8'h00;
    ff_ram[11311] = 8'h00;
    ff_ram[11312] = 8'h00;
    ff_ram[11313] = 8'h00;
    ff_ram[11314] = 8'h00;
    ff_ram[11315] = 8'h00;
    ff_ram[11316] = 8'h00;
    ff_ram[11317] = 8'h00;
    ff_ram[11318] = 8'h00;
    ff_ram[11319] = 8'h00;
    ff_ram[11320] = 8'h00;
    ff_ram[11321] = 8'h00;
    ff_ram[11322] = 8'h00;
    ff_ram[11323] = 8'h00;
    ff_ram[11324] = 8'h00;
    ff_ram[11325] = 8'h00;
    ff_ram[11326] = 8'h00;
    ff_ram[11327] = 8'h00;
    ff_ram[11328] = 8'h00;
    ff_ram[11329] = 8'h00;
    ff_ram[11330] = 8'h00;
    ff_ram[11331] = 8'h00;
    ff_ram[11332] = 8'h00;
    ff_ram[11333] = 8'h00;
    ff_ram[11334] = 8'h00;
    ff_ram[11335] = 8'h00;
    ff_ram[11336] = 8'h00;
    ff_ram[11337] = 8'h00;
    ff_ram[11338] = 8'h00;
    ff_ram[11339] = 8'h00;
    ff_ram[11340] = 8'h00;
    ff_ram[11341] = 8'h00;
    ff_ram[11342] = 8'h00;
    ff_ram[11343] = 8'h00;
    ff_ram[11344] = 8'h00;
    ff_ram[11345] = 8'h00;
    ff_ram[11346] = 8'h00;
    ff_ram[11347] = 8'h00;
    ff_ram[11348] = 8'h00;
    ff_ram[11349] = 8'h00;
    ff_ram[11350] = 8'h00;
    ff_ram[11351] = 8'h00;
    ff_ram[11352] = 8'h00;
    ff_ram[11353] = 8'h00;
    ff_ram[11354] = 8'h00;
    ff_ram[11355] = 8'h00;
    ff_ram[11356] = 8'h00;
    ff_ram[11357] = 8'h00;
    ff_ram[11358] = 8'h00;
    ff_ram[11359] = 8'h00;
    ff_ram[11360] = 8'h00;
    ff_ram[11361] = 8'h00;
    ff_ram[11362] = 8'h00;
    ff_ram[11363] = 8'h00;
    ff_ram[11364] = 8'h00;
    ff_ram[11365] = 8'h00;
    ff_ram[11366] = 8'h00;
    ff_ram[11367] = 8'h00;
    ff_ram[11368] = 8'h00;
    ff_ram[11369] = 8'h00;
    ff_ram[11370] = 8'h00;
    ff_ram[11371] = 8'h00;
    ff_ram[11372] = 8'h00;
    ff_ram[11373] = 8'h00;
    ff_ram[11374] = 8'h00;
    ff_ram[11375] = 8'h00;
    ff_ram[11376] = 8'h00;
    ff_ram[11377] = 8'h00;
    ff_ram[11378] = 8'h00;
    ff_ram[11379] = 8'h00;
    ff_ram[11380] = 8'h00;
    ff_ram[11381] = 8'h00;
    ff_ram[11382] = 8'h00;
    ff_ram[11383] = 8'h00;
    ff_ram[11384] = 8'h00;
    ff_ram[11385] = 8'h00;
    ff_ram[11386] = 8'h00;
    ff_ram[11387] = 8'h00;
    ff_ram[11388] = 8'h00;
    ff_ram[11389] = 8'h00;
    ff_ram[11390] = 8'h00;
    ff_ram[11391] = 8'h00;
    ff_ram[11392] = 8'h00;
    ff_ram[11393] = 8'h00;
    ff_ram[11394] = 8'h00;
    ff_ram[11395] = 8'h00;
    ff_ram[11396] = 8'h00;
    ff_ram[11397] = 8'h00;
    ff_ram[11398] = 8'h00;
    ff_ram[11399] = 8'h00;
    ff_ram[11400] = 8'h00;
    ff_ram[11401] = 8'h00;
    ff_ram[11402] = 8'h00;
    ff_ram[11403] = 8'h00;
    ff_ram[11404] = 8'h00;
    ff_ram[11405] = 8'h00;
    ff_ram[11406] = 8'h00;
    ff_ram[11407] = 8'h00;
    ff_ram[11408] = 8'h00;
    ff_ram[11409] = 8'h00;
    ff_ram[11410] = 8'h00;
    ff_ram[11411] = 8'h00;
    ff_ram[11412] = 8'h00;
    ff_ram[11413] = 8'h00;
    ff_ram[11414] = 8'h00;
    ff_ram[11415] = 8'h00;
    ff_ram[11416] = 8'h00;
    ff_ram[11417] = 8'h00;
    ff_ram[11418] = 8'h00;
    ff_ram[11419] = 8'h00;
    ff_ram[11420] = 8'h00;
    ff_ram[11421] = 8'h00;
    ff_ram[11422] = 8'h00;
    ff_ram[11423] = 8'h00;
    ff_ram[11424] = 8'h00;
    ff_ram[11425] = 8'h00;
    ff_ram[11426] = 8'h00;
    ff_ram[11427] = 8'h00;
    ff_ram[11428] = 8'h00;
    ff_ram[11429] = 8'h00;
    ff_ram[11430] = 8'h00;
    ff_ram[11431] = 8'h00;
    ff_ram[11432] = 8'h00;
    ff_ram[11433] = 8'h00;
    ff_ram[11434] = 8'h00;
    ff_ram[11435] = 8'h00;
    ff_ram[11436] = 8'h00;
    ff_ram[11437] = 8'h00;
    ff_ram[11438] = 8'h00;
    ff_ram[11439] = 8'h00;
    ff_ram[11440] = 8'h00;
    ff_ram[11441] = 8'h00;
    ff_ram[11442] = 8'h00;
    ff_ram[11443] = 8'h00;
    ff_ram[11444] = 8'h00;
    ff_ram[11445] = 8'h00;
    ff_ram[11446] = 8'h00;
    ff_ram[11447] = 8'h00;
    ff_ram[11448] = 8'h00;
    ff_ram[11449] = 8'h00;
    ff_ram[11450] = 8'h00;
    ff_ram[11451] = 8'h00;
    ff_ram[11452] = 8'h00;
    ff_ram[11453] = 8'h00;
    ff_ram[11454] = 8'h00;
    ff_ram[11455] = 8'h00;
    ff_ram[11456] = 8'h00;
    ff_ram[11457] = 8'h00;
    ff_ram[11458] = 8'h00;
    ff_ram[11459] = 8'h00;
    ff_ram[11460] = 8'h00;
    ff_ram[11461] = 8'h00;
    ff_ram[11462] = 8'h00;
    ff_ram[11463] = 8'h00;
    ff_ram[11464] = 8'h00;
    ff_ram[11465] = 8'h00;
    ff_ram[11466] = 8'h00;
    ff_ram[11467] = 8'h00;
    ff_ram[11468] = 8'h00;
    ff_ram[11469] = 8'h00;
    ff_ram[11470] = 8'h00;
    ff_ram[11471] = 8'h00;
    ff_ram[11472] = 8'h00;
    ff_ram[11473] = 8'h00;
    ff_ram[11474] = 8'h00;
    ff_ram[11475] = 8'h00;
    ff_ram[11476] = 8'h00;
    ff_ram[11477] = 8'h00;
    ff_ram[11478] = 8'h00;
    ff_ram[11479] = 8'h00;
    ff_ram[11480] = 8'h00;
    ff_ram[11481] = 8'h00;
    ff_ram[11482] = 8'h00;
    ff_ram[11483] = 8'h00;
    ff_ram[11484] = 8'h00;
    ff_ram[11485] = 8'h00;
    ff_ram[11486] = 8'h00;
    ff_ram[11487] = 8'h00;
    ff_ram[11488] = 8'h00;
    ff_ram[11489] = 8'h00;
    ff_ram[11490] = 8'h00;
    ff_ram[11491] = 8'h00;
    ff_ram[11492] = 8'h00;
    ff_ram[11493] = 8'h00;
    ff_ram[11494] = 8'h00;
    ff_ram[11495] = 8'h00;
    ff_ram[11496] = 8'h00;
    ff_ram[11497] = 8'h00;
    ff_ram[11498] = 8'h00;
    ff_ram[11499] = 8'h00;
    ff_ram[11500] = 8'h00;
    ff_ram[11501] = 8'h00;
    ff_ram[11502] = 8'h00;
    ff_ram[11503] = 8'h00;
    ff_ram[11504] = 8'h00;
    ff_ram[11505] = 8'h00;
    ff_ram[11506] = 8'h00;
    ff_ram[11507] = 8'h00;
    ff_ram[11508] = 8'h00;
    ff_ram[11509] = 8'h00;
    ff_ram[11510] = 8'h00;
    ff_ram[11511] = 8'h00;
    ff_ram[11512] = 8'h00;
    ff_ram[11513] = 8'h00;
    ff_ram[11514] = 8'h00;
    ff_ram[11515] = 8'h00;
    ff_ram[11516] = 8'h00;
    ff_ram[11517] = 8'h00;
    ff_ram[11518] = 8'h00;
    ff_ram[11519] = 8'h00;
    ff_ram[11520] = 8'h00;
    ff_ram[11521] = 8'h00;
    ff_ram[11522] = 8'h00;
    ff_ram[11523] = 8'h00;
    ff_ram[11524] = 8'h00;
    ff_ram[11525] = 8'h00;
    ff_ram[11526] = 8'h00;
    ff_ram[11527] = 8'h00;
    ff_ram[11528] = 8'h00;
    ff_ram[11529] = 8'h00;
    ff_ram[11530] = 8'h00;
    ff_ram[11531] = 8'h00;
    ff_ram[11532] = 8'h00;
    ff_ram[11533] = 8'h00;
    ff_ram[11534] = 8'h00;
    ff_ram[11535] = 8'h00;
    ff_ram[11536] = 8'h00;
    ff_ram[11537] = 8'h00;
    ff_ram[11538] = 8'h00;
    ff_ram[11539] = 8'h00;
    ff_ram[11540] = 8'h00;
    ff_ram[11541] = 8'h00;
    ff_ram[11542] = 8'h00;
    ff_ram[11543] = 8'h00;
    ff_ram[11544] = 8'h00;
    ff_ram[11545] = 8'h00;
    ff_ram[11546] = 8'h00;
    ff_ram[11547] = 8'h00;
    ff_ram[11548] = 8'h00;
    ff_ram[11549] = 8'h00;
    ff_ram[11550] = 8'h00;
    ff_ram[11551] = 8'h00;
    ff_ram[11552] = 8'h00;
    ff_ram[11553] = 8'h00;
    ff_ram[11554] = 8'h00;
    ff_ram[11555] = 8'h00;
    ff_ram[11556] = 8'h00;
    ff_ram[11557] = 8'h00;
    ff_ram[11558] = 8'h00;
    ff_ram[11559] = 8'h00;
    ff_ram[11560] = 8'h00;
    ff_ram[11561] = 8'h00;
    ff_ram[11562] = 8'h00;
    ff_ram[11563] = 8'h00;
    ff_ram[11564] = 8'h00;
    ff_ram[11565] = 8'h00;
    ff_ram[11566] = 8'h00;
    ff_ram[11567] = 8'h00;
    ff_ram[11568] = 8'h00;
    ff_ram[11569] = 8'h00;
    ff_ram[11570] = 8'h00;
    ff_ram[11571] = 8'h00;
    ff_ram[11572] = 8'h00;
    ff_ram[11573] = 8'h00;
    ff_ram[11574] = 8'h00;
    ff_ram[11575] = 8'h00;
    ff_ram[11576] = 8'h00;
    ff_ram[11577] = 8'h00;
    ff_ram[11578] = 8'h00;
    ff_ram[11579] = 8'h00;
    ff_ram[11580] = 8'h00;
    ff_ram[11581] = 8'h00;
    ff_ram[11582] = 8'h00;
    ff_ram[11583] = 8'h00;
    ff_ram[11584] = 8'h00;
    ff_ram[11585] = 8'h00;
    ff_ram[11586] = 8'h00;
    ff_ram[11587] = 8'h00;
    ff_ram[11588] = 8'h00;
    ff_ram[11589] = 8'h00;
    ff_ram[11590] = 8'h00;
    ff_ram[11591] = 8'h00;
    ff_ram[11592] = 8'h00;
    ff_ram[11593] = 8'h00;
    ff_ram[11594] = 8'h00;
    ff_ram[11595] = 8'h00;
    ff_ram[11596] = 8'h00;
    ff_ram[11597] = 8'h00;
    ff_ram[11598] = 8'h00;
    ff_ram[11599] = 8'h00;
    ff_ram[11600] = 8'h00;
    ff_ram[11601] = 8'h00;
    ff_ram[11602] = 8'h00;
    ff_ram[11603] = 8'h00;
    ff_ram[11604] = 8'h00;
    ff_ram[11605] = 8'h00;
    ff_ram[11606] = 8'h00;
    ff_ram[11607] = 8'h00;
    ff_ram[11608] = 8'h00;
    ff_ram[11609] = 8'h00;
    ff_ram[11610] = 8'h00;
    ff_ram[11611] = 8'h00;
    ff_ram[11612] = 8'h00;
    ff_ram[11613] = 8'h00;
    ff_ram[11614] = 8'h00;
    ff_ram[11615] = 8'h00;
    ff_ram[11616] = 8'h00;
    ff_ram[11617] = 8'h00;
    ff_ram[11618] = 8'h00;
    ff_ram[11619] = 8'h00;
    ff_ram[11620] = 8'h00;
    ff_ram[11621] = 8'h00;
    ff_ram[11622] = 8'h00;
    ff_ram[11623] = 8'h00;
    ff_ram[11624] = 8'h00;
    ff_ram[11625] = 8'h00;
    ff_ram[11626] = 8'h00;
    ff_ram[11627] = 8'h00;
    ff_ram[11628] = 8'h00;
    ff_ram[11629] = 8'h00;
    ff_ram[11630] = 8'h00;
    ff_ram[11631] = 8'h00;
    ff_ram[11632] = 8'h00;
    ff_ram[11633] = 8'h00;
    ff_ram[11634] = 8'h00;
    ff_ram[11635] = 8'h00;
    ff_ram[11636] = 8'h00;
    ff_ram[11637] = 8'h00;
    ff_ram[11638] = 8'h00;
    ff_ram[11639] = 8'h00;
    ff_ram[11640] = 8'h00;
    ff_ram[11641] = 8'h00;
    ff_ram[11642] = 8'h00;
    ff_ram[11643] = 8'h00;
    ff_ram[11644] = 8'h00;
    ff_ram[11645] = 8'h00;
    ff_ram[11646] = 8'h00;
    ff_ram[11647] = 8'h00;
    ff_ram[11648] = 8'h00;
    ff_ram[11649] = 8'h00;
    ff_ram[11650] = 8'h00;
    ff_ram[11651] = 8'h00;
    ff_ram[11652] = 8'h00;
    ff_ram[11653] = 8'h00;
    ff_ram[11654] = 8'h00;
    ff_ram[11655] = 8'h00;
    ff_ram[11656] = 8'h00;
    ff_ram[11657] = 8'h00;
    ff_ram[11658] = 8'h00;
    ff_ram[11659] = 8'h00;
    ff_ram[11660] = 8'h00;
    ff_ram[11661] = 8'h00;
    ff_ram[11662] = 8'h00;
    ff_ram[11663] = 8'h00;
    ff_ram[11664] = 8'h00;
    ff_ram[11665] = 8'h00;
    ff_ram[11666] = 8'h00;
    ff_ram[11667] = 8'h00;
    ff_ram[11668] = 8'h00;
    ff_ram[11669] = 8'h00;
    ff_ram[11670] = 8'h00;
    ff_ram[11671] = 8'h00;
    ff_ram[11672] = 8'h00;
    ff_ram[11673] = 8'h00;
    ff_ram[11674] = 8'h00;
    ff_ram[11675] = 8'h00;
    ff_ram[11676] = 8'h00;
    ff_ram[11677] = 8'h00;
    ff_ram[11678] = 8'h00;
    ff_ram[11679] = 8'h00;
    ff_ram[11680] = 8'h00;
    ff_ram[11681] = 8'h00;
    ff_ram[11682] = 8'h00;
    ff_ram[11683] = 8'h00;
    ff_ram[11684] = 8'h00;
    ff_ram[11685] = 8'h00;
    ff_ram[11686] = 8'h00;
    ff_ram[11687] = 8'h00;
    ff_ram[11688] = 8'h00;
    ff_ram[11689] = 8'h00;
    ff_ram[11690] = 8'h00;
    ff_ram[11691] = 8'h00;
    ff_ram[11692] = 8'h00;
    ff_ram[11693] = 8'h00;
    ff_ram[11694] = 8'h00;
    ff_ram[11695] = 8'h00;
    ff_ram[11696] = 8'h00;
    ff_ram[11697] = 8'h00;
    ff_ram[11698] = 8'h00;
    ff_ram[11699] = 8'h00;
    ff_ram[11700] = 8'h00;
    ff_ram[11701] = 8'h00;
    ff_ram[11702] = 8'h00;
    ff_ram[11703] = 8'h00;
    ff_ram[11704] = 8'h00;
    ff_ram[11705] = 8'h00;
    ff_ram[11706] = 8'h00;
    ff_ram[11707] = 8'h00;
    ff_ram[11708] = 8'h00;
    ff_ram[11709] = 8'h00;
    ff_ram[11710] = 8'h00;
    ff_ram[11711] = 8'h00;
    ff_ram[11712] = 8'h00;
    ff_ram[11713] = 8'h00;
    ff_ram[11714] = 8'h00;
    ff_ram[11715] = 8'h00;
    ff_ram[11716] = 8'h00;
    ff_ram[11717] = 8'h00;
    ff_ram[11718] = 8'h00;
    ff_ram[11719] = 8'h00;
    ff_ram[11720] = 8'h00;
    ff_ram[11721] = 8'h00;
    ff_ram[11722] = 8'h00;
    ff_ram[11723] = 8'h00;
    ff_ram[11724] = 8'h00;
    ff_ram[11725] = 8'h00;
    ff_ram[11726] = 8'h00;
    ff_ram[11727] = 8'h00;
    ff_ram[11728] = 8'h00;
    ff_ram[11729] = 8'h00;
    ff_ram[11730] = 8'h00;
    ff_ram[11731] = 8'h00;
    ff_ram[11732] = 8'h00;
    ff_ram[11733] = 8'h00;
    ff_ram[11734] = 8'h00;
    ff_ram[11735] = 8'h00;
    ff_ram[11736] = 8'h00;
    ff_ram[11737] = 8'h00;
    ff_ram[11738] = 8'h00;
    ff_ram[11739] = 8'h00;
    ff_ram[11740] = 8'h00;
    ff_ram[11741] = 8'h00;
    ff_ram[11742] = 8'h00;
    ff_ram[11743] = 8'h00;
    ff_ram[11744] = 8'h00;
    ff_ram[11745] = 8'h00;
    ff_ram[11746] = 8'h00;
    ff_ram[11747] = 8'h00;
    ff_ram[11748] = 8'h00;
    ff_ram[11749] = 8'h00;
    ff_ram[11750] = 8'h00;
    ff_ram[11751] = 8'h00;
    ff_ram[11752] = 8'h00;
    ff_ram[11753] = 8'h00;
    ff_ram[11754] = 8'h00;
    ff_ram[11755] = 8'h00;
    ff_ram[11756] = 8'h00;
    ff_ram[11757] = 8'h00;
    ff_ram[11758] = 8'h00;
    ff_ram[11759] = 8'h00;
    ff_ram[11760] = 8'h00;
    ff_ram[11761] = 8'h00;
    ff_ram[11762] = 8'h00;
    ff_ram[11763] = 8'h00;
    ff_ram[11764] = 8'h00;
    ff_ram[11765] = 8'h00;
    ff_ram[11766] = 8'h00;
    ff_ram[11767] = 8'h00;
    ff_ram[11768] = 8'h00;
    ff_ram[11769] = 8'h00;
    ff_ram[11770] = 8'h00;
    ff_ram[11771] = 8'h00;
    ff_ram[11772] = 8'h00;
    ff_ram[11773] = 8'h00;
    ff_ram[11774] = 8'h00;
    ff_ram[11775] = 8'h00;
    ff_ram[11776] = 8'h00;
    ff_ram[11777] = 8'h00;
    ff_ram[11778] = 8'h00;
    ff_ram[11779] = 8'h00;
    ff_ram[11780] = 8'h00;
    ff_ram[11781] = 8'h00;
    ff_ram[11782] = 8'h00;
    ff_ram[11783] = 8'h00;
    ff_ram[11784] = 8'h00;
    ff_ram[11785] = 8'h00;
    ff_ram[11786] = 8'h00;
    ff_ram[11787] = 8'h00;
    ff_ram[11788] = 8'h00;
    ff_ram[11789] = 8'h00;
    ff_ram[11790] = 8'h00;
    ff_ram[11791] = 8'h00;
    ff_ram[11792] = 8'h00;
    ff_ram[11793] = 8'h00;
    ff_ram[11794] = 8'h00;
    ff_ram[11795] = 8'h00;
    ff_ram[11796] = 8'h00;
    ff_ram[11797] = 8'h00;
    ff_ram[11798] = 8'h00;
    ff_ram[11799] = 8'h00;
    ff_ram[11800] = 8'h00;
    ff_ram[11801] = 8'h00;
    ff_ram[11802] = 8'h00;
    ff_ram[11803] = 8'h00;
    ff_ram[11804] = 8'h00;
    ff_ram[11805] = 8'h00;
    ff_ram[11806] = 8'h00;
    ff_ram[11807] = 8'h00;
    ff_ram[11808] = 8'h00;
    ff_ram[11809] = 8'h00;
    ff_ram[11810] = 8'h00;
    ff_ram[11811] = 8'h00;
    ff_ram[11812] = 8'h00;
    ff_ram[11813] = 8'h00;
    ff_ram[11814] = 8'h00;
    ff_ram[11815] = 8'h00;
    ff_ram[11816] = 8'h00;
    ff_ram[11817] = 8'h00;
    ff_ram[11818] = 8'h00;
    ff_ram[11819] = 8'h00;
    ff_ram[11820] = 8'h00;
    ff_ram[11821] = 8'h00;
    ff_ram[11822] = 8'h00;
    ff_ram[11823] = 8'h00;
    ff_ram[11824] = 8'h00;
    ff_ram[11825] = 8'h00;
    ff_ram[11826] = 8'h00;
    ff_ram[11827] = 8'h00;
    ff_ram[11828] = 8'h00;
    ff_ram[11829] = 8'h00;
    ff_ram[11830] = 8'h00;
    ff_ram[11831] = 8'h00;
    ff_ram[11832] = 8'h00;
    ff_ram[11833] = 8'h00;
    ff_ram[11834] = 8'h00;
    ff_ram[11835] = 8'h00;
    ff_ram[11836] = 8'h00;
    ff_ram[11837] = 8'h00;
    ff_ram[11838] = 8'h00;
    ff_ram[11839] = 8'h00;
    ff_ram[11840] = 8'h00;
    ff_ram[11841] = 8'h00;
    ff_ram[11842] = 8'h00;
    ff_ram[11843] = 8'h00;
    ff_ram[11844] = 8'h00;
    ff_ram[11845] = 8'h00;
    ff_ram[11846] = 8'h00;
    ff_ram[11847] = 8'h00;
    ff_ram[11848] = 8'h00;
    ff_ram[11849] = 8'h00;
    ff_ram[11850] = 8'h00;
    ff_ram[11851] = 8'h00;
    ff_ram[11852] = 8'h00;
    ff_ram[11853] = 8'h00;
    ff_ram[11854] = 8'h00;
    ff_ram[11855] = 8'h00;
    ff_ram[11856] = 8'h00;
    ff_ram[11857] = 8'h00;
    ff_ram[11858] = 8'h00;
    ff_ram[11859] = 8'h00;
    ff_ram[11860] = 8'h00;
    ff_ram[11861] = 8'h00;
    ff_ram[11862] = 8'h00;
    ff_ram[11863] = 8'h00;
    ff_ram[11864] = 8'h00;
    ff_ram[11865] = 8'h00;
    ff_ram[11866] = 8'h00;
    ff_ram[11867] = 8'h00;
    ff_ram[11868] = 8'h00;
    ff_ram[11869] = 8'h00;
    ff_ram[11870] = 8'h00;
    ff_ram[11871] = 8'h00;
    ff_ram[11872] = 8'h00;
    ff_ram[11873] = 8'h00;
    ff_ram[11874] = 8'h00;
    ff_ram[11875] = 8'h00;
    ff_ram[11876] = 8'h00;
    ff_ram[11877] = 8'h00;
    ff_ram[11878] = 8'h00;
    ff_ram[11879] = 8'h00;
    ff_ram[11880] = 8'h00;
    ff_ram[11881] = 8'h00;
    ff_ram[11882] = 8'h00;
    ff_ram[11883] = 8'h00;
    ff_ram[11884] = 8'h00;
    ff_ram[11885] = 8'h00;
    ff_ram[11886] = 8'h00;
    ff_ram[11887] = 8'h00;
    ff_ram[11888] = 8'h00;
    ff_ram[11889] = 8'h00;
    ff_ram[11890] = 8'h00;
    ff_ram[11891] = 8'h00;
    ff_ram[11892] = 8'h00;
    ff_ram[11893] = 8'h00;
    ff_ram[11894] = 8'h00;
    ff_ram[11895] = 8'h00;
    ff_ram[11896] = 8'h00;
    ff_ram[11897] = 8'h00;
    ff_ram[11898] = 8'h00;
    ff_ram[11899] = 8'h00;
    ff_ram[11900] = 8'h00;
    ff_ram[11901] = 8'h00;
    ff_ram[11902] = 8'h00;
    ff_ram[11903] = 8'h00;
    ff_ram[11904] = 8'h00;
    ff_ram[11905] = 8'h00;
    ff_ram[11906] = 8'h00;
    ff_ram[11907] = 8'h00;
    ff_ram[11908] = 8'h00;
    ff_ram[11909] = 8'h00;
    ff_ram[11910] = 8'h00;
    ff_ram[11911] = 8'h00;
    ff_ram[11912] = 8'h00;
    ff_ram[11913] = 8'h00;
    ff_ram[11914] = 8'h00;
    ff_ram[11915] = 8'h00;
    ff_ram[11916] = 8'h00;
    ff_ram[11917] = 8'h00;
    ff_ram[11918] = 8'h00;
    ff_ram[11919] = 8'h00;
    ff_ram[11920] = 8'h00;
    ff_ram[11921] = 8'h00;
    ff_ram[11922] = 8'h00;
    ff_ram[11923] = 8'h00;
    ff_ram[11924] = 8'h00;
    ff_ram[11925] = 8'h00;
    ff_ram[11926] = 8'h00;
    ff_ram[11927] = 8'h00;
    ff_ram[11928] = 8'h00;
    ff_ram[11929] = 8'h00;
    ff_ram[11930] = 8'h00;
    ff_ram[11931] = 8'h00;
    ff_ram[11932] = 8'h00;
    ff_ram[11933] = 8'h00;
    ff_ram[11934] = 8'h00;
    ff_ram[11935] = 8'h00;
    ff_ram[11936] = 8'h00;
    ff_ram[11937] = 8'h00;
    ff_ram[11938] = 8'h00;
    ff_ram[11939] = 8'h00;
    ff_ram[11940] = 8'h00;
    ff_ram[11941] = 8'h00;
    ff_ram[11942] = 8'h00;
    ff_ram[11943] = 8'h00;
    ff_ram[11944] = 8'h00;
    ff_ram[11945] = 8'h00;
    ff_ram[11946] = 8'h00;
    ff_ram[11947] = 8'h00;
    ff_ram[11948] = 8'h00;
    ff_ram[11949] = 8'h00;
    ff_ram[11950] = 8'h00;
    ff_ram[11951] = 8'h00;
    ff_ram[11952] = 8'h00;
    ff_ram[11953] = 8'h00;
    ff_ram[11954] = 8'h00;
    ff_ram[11955] = 8'h00;
    ff_ram[11956] = 8'h00;
    ff_ram[11957] = 8'h00;
    ff_ram[11958] = 8'h00;
    ff_ram[11959] = 8'h00;
    ff_ram[11960] = 8'h00;
    ff_ram[11961] = 8'h00;
    ff_ram[11962] = 8'h00;
    ff_ram[11963] = 8'h00;
    ff_ram[11964] = 8'h00;
    ff_ram[11965] = 8'h00;
    ff_ram[11966] = 8'h00;
    ff_ram[11967] = 8'h00;
    ff_ram[11968] = 8'h00;
    ff_ram[11969] = 8'h00;
    ff_ram[11970] = 8'h00;
    ff_ram[11971] = 8'h00;
    ff_ram[11972] = 8'h00;
    ff_ram[11973] = 8'h00;
    ff_ram[11974] = 8'h00;
    ff_ram[11975] = 8'h00;
    ff_ram[11976] = 8'h00;
    ff_ram[11977] = 8'h00;
    ff_ram[11978] = 8'h00;
    ff_ram[11979] = 8'h00;
    ff_ram[11980] = 8'h00;
    ff_ram[11981] = 8'h00;
    ff_ram[11982] = 8'h00;
    ff_ram[11983] = 8'h00;
    ff_ram[11984] = 8'h00;
    ff_ram[11985] = 8'h00;
    ff_ram[11986] = 8'h00;
    ff_ram[11987] = 8'h00;
    ff_ram[11988] = 8'h00;
    ff_ram[11989] = 8'h00;
    ff_ram[11990] = 8'h00;
    ff_ram[11991] = 8'h00;
    ff_ram[11992] = 8'h00;
    ff_ram[11993] = 8'h00;
    ff_ram[11994] = 8'h00;
    ff_ram[11995] = 8'h00;
    ff_ram[11996] = 8'h00;
    ff_ram[11997] = 8'h00;
    ff_ram[11998] = 8'h00;
    ff_ram[11999] = 8'h00;
    ff_ram[12000] = 8'h00;
    ff_ram[12001] = 8'h00;
    ff_ram[12002] = 8'h00;
    ff_ram[12003] = 8'h00;
    ff_ram[12004] = 8'h00;
    ff_ram[12005] = 8'h00;
    ff_ram[12006] = 8'h00;
    ff_ram[12007] = 8'h00;
    ff_ram[12008] = 8'h00;
    ff_ram[12009] = 8'h00;
    ff_ram[12010] = 8'h00;
    ff_ram[12011] = 8'h00;
    ff_ram[12012] = 8'h00;
    ff_ram[12013] = 8'h00;
    ff_ram[12014] = 8'h00;
    ff_ram[12015] = 8'h00;
    ff_ram[12016] = 8'h00;
    ff_ram[12017] = 8'h00;
    ff_ram[12018] = 8'h00;
    ff_ram[12019] = 8'h00;
    ff_ram[12020] = 8'h00;
    ff_ram[12021] = 8'h00;
    ff_ram[12022] = 8'h00;
    ff_ram[12023] = 8'h00;
    ff_ram[12024] = 8'h00;
    ff_ram[12025] = 8'h00;
    ff_ram[12026] = 8'h00;
    ff_ram[12027] = 8'h00;
    ff_ram[12028] = 8'h00;
    ff_ram[12029] = 8'h00;
    ff_ram[12030] = 8'h00;
    ff_ram[12031] = 8'h00;
    ff_ram[12032] = 8'h00;
    ff_ram[12033] = 8'h00;
    ff_ram[12034] = 8'h00;
    ff_ram[12035] = 8'h00;
    ff_ram[12036] = 8'h00;
    ff_ram[12037] = 8'h00;
    ff_ram[12038] = 8'h00;
    ff_ram[12039] = 8'h00;
    ff_ram[12040] = 8'h00;
    ff_ram[12041] = 8'h00;
    ff_ram[12042] = 8'h00;
    ff_ram[12043] = 8'h00;
    ff_ram[12044] = 8'h00;
    ff_ram[12045] = 8'h00;
    ff_ram[12046] = 8'h00;
    ff_ram[12047] = 8'h00;
    ff_ram[12048] = 8'h00;
    ff_ram[12049] = 8'h00;
    ff_ram[12050] = 8'h00;
    ff_ram[12051] = 8'h00;
    ff_ram[12052] = 8'h00;
    ff_ram[12053] = 8'h00;
    ff_ram[12054] = 8'h00;
    ff_ram[12055] = 8'h00;
    ff_ram[12056] = 8'h00;
    ff_ram[12057] = 8'h00;
    ff_ram[12058] = 8'h00;
    ff_ram[12059] = 8'h00;
    ff_ram[12060] = 8'h00;
    ff_ram[12061] = 8'h00;
    ff_ram[12062] = 8'h00;
    ff_ram[12063] = 8'h00;
    ff_ram[12064] = 8'h00;
    ff_ram[12065] = 8'h00;
    ff_ram[12066] = 8'h00;
    ff_ram[12067] = 8'h00;
    ff_ram[12068] = 8'h00;
    ff_ram[12069] = 8'h00;
    ff_ram[12070] = 8'h00;
    ff_ram[12071] = 8'h00;
    ff_ram[12072] = 8'h00;
    ff_ram[12073] = 8'h00;
    ff_ram[12074] = 8'h00;
    ff_ram[12075] = 8'h00;
    ff_ram[12076] = 8'h00;
    ff_ram[12077] = 8'h00;
    ff_ram[12078] = 8'h00;
    ff_ram[12079] = 8'h00;
    ff_ram[12080] = 8'h00;
    ff_ram[12081] = 8'h00;
    ff_ram[12082] = 8'h00;
    ff_ram[12083] = 8'h00;
    ff_ram[12084] = 8'h00;
    ff_ram[12085] = 8'h00;
    ff_ram[12086] = 8'h00;
    ff_ram[12087] = 8'h00;
    ff_ram[12088] = 8'h00;
    ff_ram[12089] = 8'h00;
    ff_ram[12090] = 8'h00;
    ff_ram[12091] = 8'h00;
    ff_ram[12092] = 8'h00;
    ff_ram[12093] = 8'h00;
    ff_ram[12094] = 8'h00;
    ff_ram[12095] = 8'h00;
    ff_ram[12096] = 8'h00;
    ff_ram[12097] = 8'h00;
    ff_ram[12098] = 8'h00;
    ff_ram[12099] = 8'h00;
    ff_ram[12100] = 8'h00;
    ff_ram[12101] = 8'h00;
    ff_ram[12102] = 8'h00;
    ff_ram[12103] = 8'h00;
    ff_ram[12104] = 8'h00;
    ff_ram[12105] = 8'h00;
    ff_ram[12106] = 8'h00;
    ff_ram[12107] = 8'h00;
    ff_ram[12108] = 8'h00;
    ff_ram[12109] = 8'h00;
    ff_ram[12110] = 8'h00;
    ff_ram[12111] = 8'h00;
    ff_ram[12112] = 8'h00;
    ff_ram[12113] = 8'h00;
    ff_ram[12114] = 8'h00;
    ff_ram[12115] = 8'h00;
    ff_ram[12116] = 8'h00;
    ff_ram[12117] = 8'h00;
    ff_ram[12118] = 8'h00;
    ff_ram[12119] = 8'h00;
    ff_ram[12120] = 8'h00;
    ff_ram[12121] = 8'h00;
    ff_ram[12122] = 8'h00;
    ff_ram[12123] = 8'h00;
    ff_ram[12124] = 8'h00;
    ff_ram[12125] = 8'h00;
    ff_ram[12126] = 8'h00;
    ff_ram[12127] = 8'h00;
    ff_ram[12128] = 8'h00;
    ff_ram[12129] = 8'h00;
    ff_ram[12130] = 8'h00;
    ff_ram[12131] = 8'h00;
    ff_ram[12132] = 8'h00;
    ff_ram[12133] = 8'h00;
    ff_ram[12134] = 8'h00;
    ff_ram[12135] = 8'h00;
    ff_ram[12136] = 8'h00;
    ff_ram[12137] = 8'h00;
    ff_ram[12138] = 8'h00;
    ff_ram[12139] = 8'h00;
    ff_ram[12140] = 8'h00;
    ff_ram[12141] = 8'h00;
    ff_ram[12142] = 8'h00;
    ff_ram[12143] = 8'h00;
    ff_ram[12144] = 8'h00;
    ff_ram[12145] = 8'h00;
    ff_ram[12146] = 8'h00;
    ff_ram[12147] = 8'h00;
    ff_ram[12148] = 8'h00;
    ff_ram[12149] = 8'h00;
    ff_ram[12150] = 8'h00;
    ff_ram[12151] = 8'h00;
    ff_ram[12152] = 8'h00;
    ff_ram[12153] = 8'h00;
    ff_ram[12154] = 8'h00;
    ff_ram[12155] = 8'h00;
    ff_ram[12156] = 8'h00;
    ff_ram[12157] = 8'h00;
    ff_ram[12158] = 8'h00;
    ff_ram[12159] = 8'h00;
    ff_ram[12160] = 8'h00;
    ff_ram[12161] = 8'h00;
    ff_ram[12162] = 8'h00;
    ff_ram[12163] = 8'h00;
    ff_ram[12164] = 8'h00;
    ff_ram[12165] = 8'h00;
    ff_ram[12166] = 8'h00;
    ff_ram[12167] = 8'h00;
    ff_ram[12168] = 8'h00;
    ff_ram[12169] = 8'h00;
    ff_ram[12170] = 8'h00;
    ff_ram[12171] = 8'h00;
    ff_ram[12172] = 8'h00;
    ff_ram[12173] = 8'h00;
    ff_ram[12174] = 8'h00;
    ff_ram[12175] = 8'h00;
    ff_ram[12176] = 8'h00;
    ff_ram[12177] = 8'h00;
    ff_ram[12178] = 8'h00;
    ff_ram[12179] = 8'h00;
    ff_ram[12180] = 8'h00;
    ff_ram[12181] = 8'h00;
    ff_ram[12182] = 8'h00;
    ff_ram[12183] = 8'h00;
    ff_ram[12184] = 8'h00;
    ff_ram[12185] = 8'h00;
    ff_ram[12186] = 8'h00;
    ff_ram[12187] = 8'h00;
    ff_ram[12188] = 8'h00;
    ff_ram[12189] = 8'h00;
    ff_ram[12190] = 8'h00;
    ff_ram[12191] = 8'h00;
    ff_ram[12192] = 8'h00;
    ff_ram[12193] = 8'h00;
    ff_ram[12194] = 8'h00;
    ff_ram[12195] = 8'h00;
    ff_ram[12196] = 8'h00;
    ff_ram[12197] = 8'h00;
    ff_ram[12198] = 8'h00;
    ff_ram[12199] = 8'h00;
    ff_ram[12200] = 8'h00;
    ff_ram[12201] = 8'h00;
    ff_ram[12202] = 8'h00;
    ff_ram[12203] = 8'h00;
    ff_ram[12204] = 8'h00;
    ff_ram[12205] = 8'h00;
    ff_ram[12206] = 8'h00;
    ff_ram[12207] = 8'h00;
    ff_ram[12208] = 8'h00;
    ff_ram[12209] = 8'h00;
    ff_ram[12210] = 8'h00;
    ff_ram[12211] = 8'h00;
    ff_ram[12212] = 8'h00;
    ff_ram[12213] = 8'h00;
    ff_ram[12214] = 8'h00;
    ff_ram[12215] = 8'h00;
    ff_ram[12216] = 8'h00;
    ff_ram[12217] = 8'h00;
    ff_ram[12218] = 8'h00;
    ff_ram[12219] = 8'h00;
    ff_ram[12220] = 8'h00;
    ff_ram[12221] = 8'h00;
    ff_ram[12222] = 8'h00;
    ff_ram[12223] = 8'h00;
    ff_ram[12224] = 8'h00;
    ff_ram[12225] = 8'h00;
    ff_ram[12226] = 8'h00;
    ff_ram[12227] = 8'h00;
    ff_ram[12228] = 8'h00;
    ff_ram[12229] = 8'h00;
    ff_ram[12230] = 8'h00;
    ff_ram[12231] = 8'h00;
    ff_ram[12232] = 8'h00;
    ff_ram[12233] = 8'h00;
    ff_ram[12234] = 8'h00;
    ff_ram[12235] = 8'h00;
    ff_ram[12236] = 8'h00;
    ff_ram[12237] = 8'h00;
    ff_ram[12238] = 8'h00;
    ff_ram[12239] = 8'h00;
    ff_ram[12240] = 8'h00;
    ff_ram[12241] = 8'h00;
    ff_ram[12242] = 8'h00;
    ff_ram[12243] = 8'h00;
    ff_ram[12244] = 8'h00;
    ff_ram[12245] = 8'h00;
    ff_ram[12246] = 8'h00;
    ff_ram[12247] = 8'h00;
    ff_ram[12248] = 8'h00;
    ff_ram[12249] = 8'h00;
    ff_ram[12250] = 8'h00;
    ff_ram[12251] = 8'h00;
    ff_ram[12252] = 8'h00;
    ff_ram[12253] = 8'h00;
    ff_ram[12254] = 8'h00;
    ff_ram[12255] = 8'h00;
    ff_ram[12256] = 8'h00;
    ff_ram[12257] = 8'h00;
    ff_ram[12258] = 8'h00;
    ff_ram[12259] = 8'h00;
    ff_ram[12260] = 8'h00;
    ff_ram[12261] = 8'h00;
    ff_ram[12262] = 8'h00;
    ff_ram[12263] = 8'h00;
    ff_ram[12264] = 8'h00;
    ff_ram[12265] = 8'h00;
    ff_ram[12266] = 8'h00;
    ff_ram[12267] = 8'h00;
    ff_ram[12268] = 8'h00;
    ff_ram[12269] = 8'h00;
    ff_ram[12270] = 8'h00;
    ff_ram[12271] = 8'h00;
    ff_ram[12272] = 8'h00;
    ff_ram[12273] = 8'h00;
    ff_ram[12274] = 8'h00;
    ff_ram[12275] = 8'h00;
    ff_ram[12276] = 8'h00;
    ff_ram[12277] = 8'h00;
    ff_ram[12278] = 8'h00;
    ff_ram[12279] = 8'h00;
    ff_ram[12280] = 8'h00;
    ff_ram[12281] = 8'h00;
    ff_ram[12282] = 8'h00;
    ff_ram[12283] = 8'h00;
    ff_ram[12284] = 8'h00;
    ff_ram[12285] = 8'h00;
    ff_ram[12286] = 8'h00;
    ff_ram[12287] = 8'h00;
    ff_ram[12288] = 8'h00;
    ff_ram[12289] = 8'h00;
    ff_ram[12290] = 8'h00;
    ff_ram[12291] = 8'h00;
    ff_ram[12292] = 8'h00;
    ff_ram[12293] = 8'h00;
    ff_ram[12294] = 8'h00;
    ff_ram[12295] = 8'h00;
    ff_ram[12296] = 8'h00;
    ff_ram[12297] = 8'h00;
    ff_ram[12298] = 8'h00;
    ff_ram[12299] = 8'h00;
    ff_ram[12300] = 8'h00;
    ff_ram[12301] = 8'h00;
    ff_ram[12302] = 8'h00;
    ff_ram[12303] = 8'h00;
    ff_ram[12304] = 8'h00;
    ff_ram[12305] = 8'h00;
    ff_ram[12306] = 8'h00;
    ff_ram[12307] = 8'h00;
    ff_ram[12308] = 8'h00;
    ff_ram[12309] = 8'h00;
    ff_ram[12310] = 8'h00;
    ff_ram[12311] = 8'h00;
    ff_ram[12312] = 8'h00;
    ff_ram[12313] = 8'h00;
    ff_ram[12314] = 8'h00;
    ff_ram[12315] = 8'h00;
    ff_ram[12316] = 8'h00;
    ff_ram[12317] = 8'h00;
    ff_ram[12318] = 8'h00;
    ff_ram[12319] = 8'h00;
    ff_ram[12320] = 8'h00;
    ff_ram[12321] = 8'h00;
    ff_ram[12322] = 8'h00;
    ff_ram[12323] = 8'h00;
    ff_ram[12324] = 8'h00;
    ff_ram[12325] = 8'h00;
    ff_ram[12326] = 8'h00;
    ff_ram[12327] = 8'h00;
    ff_ram[12328] = 8'h00;
    ff_ram[12329] = 8'h00;
    ff_ram[12330] = 8'h00;
    ff_ram[12331] = 8'h00;
    ff_ram[12332] = 8'h00;
    ff_ram[12333] = 8'h00;
    ff_ram[12334] = 8'h00;
    ff_ram[12335] = 8'h00;
    ff_ram[12336] = 8'h00;
    ff_ram[12337] = 8'h00;
    ff_ram[12338] = 8'h00;
    ff_ram[12339] = 8'h00;
    ff_ram[12340] = 8'h00;
    ff_ram[12341] = 8'h00;
    ff_ram[12342] = 8'h00;
    ff_ram[12343] = 8'h00;
    ff_ram[12344] = 8'h00;
    ff_ram[12345] = 8'h00;
    ff_ram[12346] = 8'h00;
    ff_ram[12347] = 8'h00;
    ff_ram[12348] = 8'h00;
    ff_ram[12349] = 8'h00;
    ff_ram[12350] = 8'h00;
    ff_ram[12351] = 8'h00;
    ff_ram[12352] = 8'h00;
    ff_ram[12353] = 8'h00;
    ff_ram[12354] = 8'h00;
    ff_ram[12355] = 8'h00;
    ff_ram[12356] = 8'h00;
    ff_ram[12357] = 8'h00;
    ff_ram[12358] = 8'h00;
    ff_ram[12359] = 8'h00;
    ff_ram[12360] = 8'h00;
    ff_ram[12361] = 8'h00;
    ff_ram[12362] = 8'h00;
    ff_ram[12363] = 8'h00;
    ff_ram[12364] = 8'h00;
    ff_ram[12365] = 8'h00;
    ff_ram[12366] = 8'h00;
    ff_ram[12367] = 8'h00;
    ff_ram[12368] = 8'h00;
    ff_ram[12369] = 8'h00;
    ff_ram[12370] = 8'h00;
    ff_ram[12371] = 8'h00;
    ff_ram[12372] = 8'h00;
    ff_ram[12373] = 8'h00;
    ff_ram[12374] = 8'h00;
    ff_ram[12375] = 8'h00;
    ff_ram[12376] = 8'h00;
    ff_ram[12377] = 8'h00;
    ff_ram[12378] = 8'h00;
    ff_ram[12379] = 8'h00;
    ff_ram[12380] = 8'h00;
    ff_ram[12381] = 8'h00;
    ff_ram[12382] = 8'h00;
    ff_ram[12383] = 8'h00;
    ff_ram[12384] = 8'h00;
    ff_ram[12385] = 8'h00;
    ff_ram[12386] = 8'h00;
    ff_ram[12387] = 8'h00;
    ff_ram[12388] = 8'h00;
    ff_ram[12389] = 8'h00;
    ff_ram[12390] = 8'h00;
    ff_ram[12391] = 8'h00;
    ff_ram[12392] = 8'h00;
    ff_ram[12393] = 8'h00;
    ff_ram[12394] = 8'h00;
    ff_ram[12395] = 8'h00;
    ff_ram[12396] = 8'h00;
    ff_ram[12397] = 8'h00;
    ff_ram[12398] = 8'h00;
    ff_ram[12399] = 8'h00;
    ff_ram[12400] = 8'h00;
    ff_ram[12401] = 8'h00;
    ff_ram[12402] = 8'h00;
    ff_ram[12403] = 8'h00;
    ff_ram[12404] = 8'h00;
    ff_ram[12405] = 8'h00;
    ff_ram[12406] = 8'h00;
    ff_ram[12407] = 8'h00;
    ff_ram[12408] = 8'h00;
    ff_ram[12409] = 8'h00;
    ff_ram[12410] = 8'h00;
    ff_ram[12411] = 8'h00;
    ff_ram[12412] = 8'h00;
    ff_ram[12413] = 8'h00;
    ff_ram[12414] = 8'h00;
    ff_ram[12415] = 8'h00;
    ff_ram[12416] = 8'h00;
    ff_ram[12417] = 8'h00;
    ff_ram[12418] = 8'h00;
    ff_ram[12419] = 8'h00;
    ff_ram[12420] = 8'h00;
    ff_ram[12421] = 8'h00;
    ff_ram[12422] = 8'h00;
    ff_ram[12423] = 8'h00;
    ff_ram[12424] = 8'h00;
    ff_ram[12425] = 8'h00;
    ff_ram[12426] = 8'h00;
    ff_ram[12427] = 8'h00;
    ff_ram[12428] = 8'h00;
    ff_ram[12429] = 8'h00;
    ff_ram[12430] = 8'h00;
    ff_ram[12431] = 8'h00;
    ff_ram[12432] = 8'h00;
    ff_ram[12433] = 8'h00;
    ff_ram[12434] = 8'h00;
    ff_ram[12435] = 8'h00;
    ff_ram[12436] = 8'h00;
    ff_ram[12437] = 8'h00;
    ff_ram[12438] = 8'h00;
    ff_ram[12439] = 8'h00;
    ff_ram[12440] = 8'h00;
    ff_ram[12441] = 8'h00;
    ff_ram[12442] = 8'h00;
    ff_ram[12443] = 8'h00;
    ff_ram[12444] = 8'h00;
    ff_ram[12445] = 8'h00;
    ff_ram[12446] = 8'h00;
    ff_ram[12447] = 8'h00;
    ff_ram[12448] = 8'h00;
    ff_ram[12449] = 8'h00;
    ff_ram[12450] = 8'h00;
    ff_ram[12451] = 8'h00;
    ff_ram[12452] = 8'h00;
    ff_ram[12453] = 8'h00;
    ff_ram[12454] = 8'h00;
    ff_ram[12455] = 8'h00;
    ff_ram[12456] = 8'h00;
    ff_ram[12457] = 8'h00;
    ff_ram[12458] = 8'h00;
    ff_ram[12459] = 8'h00;
    ff_ram[12460] = 8'h00;
    ff_ram[12461] = 8'h00;
    ff_ram[12462] = 8'h00;
    ff_ram[12463] = 8'h00;
    ff_ram[12464] = 8'h00;
    ff_ram[12465] = 8'h00;
    ff_ram[12466] = 8'h00;
    ff_ram[12467] = 8'h00;
    ff_ram[12468] = 8'h00;
    ff_ram[12469] = 8'h00;
    ff_ram[12470] = 8'h00;
    ff_ram[12471] = 8'h00;
    ff_ram[12472] = 8'h00;
    ff_ram[12473] = 8'h00;
    ff_ram[12474] = 8'h00;
    ff_ram[12475] = 8'h00;
    ff_ram[12476] = 8'h00;
    ff_ram[12477] = 8'h00;
    ff_ram[12478] = 8'h00;
    ff_ram[12479] = 8'h00;
    ff_ram[12480] = 8'h00;
    ff_ram[12481] = 8'h00;
    ff_ram[12482] = 8'h00;
    ff_ram[12483] = 8'h00;
    ff_ram[12484] = 8'h00;
    ff_ram[12485] = 8'h00;
    ff_ram[12486] = 8'h00;
    ff_ram[12487] = 8'h00;
    ff_ram[12488] = 8'h00;
    ff_ram[12489] = 8'h00;
    ff_ram[12490] = 8'h00;
    ff_ram[12491] = 8'h00;
    ff_ram[12492] = 8'h00;
    ff_ram[12493] = 8'h00;
    ff_ram[12494] = 8'h00;
    ff_ram[12495] = 8'h00;
    ff_ram[12496] = 8'h00;
    ff_ram[12497] = 8'h00;
    ff_ram[12498] = 8'h00;
    ff_ram[12499] = 8'h00;
    ff_ram[12500] = 8'h00;
    ff_ram[12501] = 8'h00;
    ff_ram[12502] = 8'h00;
    ff_ram[12503] = 8'h00;
    ff_ram[12504] = 8'h00;
    ff_ram[12505] = 8'h00;
    ff_ram[12506] = 8'h00;
    ff_ram[12507] = 8'h00;
    ff_ram[12508] = 8'h00;
    ff_ram[12509] = 8'h00;
    ff_ram[12510] = 8'h00;
    ff_ram[12511] = 8'h00;
    ff_ram[12512] = 8'h00;
    ff_ram[12513] = 8'h00;
    ff_ram[12514] = 8'h00;
    ff_ram[12515] = 8'h00;
    ff_ram[12516] = 8'h00;
    ff_ram[12517] = 8'h00;
    ff_ram[12518] = 8'h00;
    ff_ram[12519] = 8'h00;
    ff_ram[12520] = 8'h00;
    ff_ram[12521] = 8'h00;
    ff_ram[12522] = 8'h00;
    ff_ram[12523] = 8'h00;
    ff_ram[12524] = 8'h00;
    ff_ram[12525] = 8'h00;
    ff_ram[12526] = 8'h00;
    ff_ram[12527] = 8'h00;
    ff_ram[12528] = 8'h00;
    ff_ram[12529] = 8'h00;
    ff_ram[12530] = 8'h00;
    ff_ram[12531] = 8'h00;
    ff_ram[12532] = 8'h00;
    ff_ram[12533] = 8'h00;
    ff_ram[12534] = 8'h00;
    ff_ram[12535] = 8'h00;
    ff_ram[12536] = 8'h00;
    ff_ram[12537] = 8'h00;
    ff_ram[12538] = 8'h00;
    ff_ram[12539] = 8'h00;
    ff_ram[12540] = 8'h00;
    ff_ram[12541] = 8'h00;
    ff_ram[12542] = 8'h00;
    ff_ram[12543] = 8'h00;
    ff_ram[12544] = 8'h00;
    ff_ram[12545] = 8'h00;
    ff_ram[12546] = 8'h00;
    ff_ram[12547] = 8'h00;
    ff_ram[12548] = 8'h00;
    ff_ram[12549] = 8'h00;
    ff_ram[12550] = 8'h00;
    ff_ram[12551] = 8'h00;
    ff_ram[12552] = 8'h00;
    ff_ram[12553] = 8'h00;
    ff_ram[12554] = 8'h00;
    ff_ram[12555] = 8'h00;
    ff_ram[12556] = 8'h00;
    ff_ram[12557] = 8'h00;
    ff_ram[12558] = 8'h00;
    ff_ram[12559] = 8'h00;
    ff_ram[12560] = 8'h00;
    ff_ram[12561] = 8'h00;
    ff_ram[12562] = 8'h00;
    ff_ram[12563] = 8'h00;
    ff_ram[12564] = 8'h00;
    ff_ram[12565] = 8'h00;
    ff_ram[12566] = 8'h00;
    ff_ram[12567] = 8'h00;
    ff_ram[12568] = 8'h00;
    ff_ram[12569] = 8'h00;
    ff_ram[12570] = 8'h00;
    ff_ram[12571] = 8'h00;
    ff_ram[12572] = 8'h00;
    ff_ram[12573] = 8'h00;
    ff_ram[12574] = 8'h00;
    ff_ram[12575] = 8'h00;
    ff_ram[12576] = 8'h00;
    ff_ram[12577] = 8'h00;
    ff_ram[12578] = 8'h00;
    ff_ram[12579] = 8'h00;
    ff_ram[12580] = 8'h00;
    ff_ram[12581] = 8'h00;
    ff_ram[12582] = 8'h00;
    ff_ram[12583] = 8'h00;
    ff_ram[12584] = 8'h00;
    ff_ram[12585] = 8'h00;
    ff_ram[12586] = 8'h00;
    ff_ram[12587] = 8'h00;
    ff_ram[12588] = 8'h00;
    ff_ram[12589] = 8'h00;
    ff_ram[12590] = 8'h00;
    ff_ram[12591] = 8'h00;
    ff_ram[12592] = 8'h00;
    ff_ram[12593] = 8'h00;
    ff_ram[12594] = 8'h00;
    ff_ram[12595] = 8'h00;
    ff_ram[12596] = 8'h00;
    ff_ram[12597] = 8'h00;
    ff_ram[12598] = 8'h00;
    ff_ram[12599] = 8'h00;
    ff_ram[12600] = 8'h00;
    ff_ram[12601] = 8'h00;
    ff_ram[12602] = 8'h00;
    ff_ram[12603] = 8'h00;
    ff_ram[12604] = 8'h00;
    ff_ram[12605] = 8'h00;
    ff_ram[12606] = 8'h00;
    ff_ram[12607] = 8'h00;
    ff_ram[12608] = 8'h00;
    ff_ram[12609] = 8'h00;
    ff_ram[12610] = 8'h00;
    ff_ram[12611] = 8'h00;
    ff_ram[12612] = 8'h00;
    ff_ram[12613] = 8'h00;
    ff_ram[12614] = 8'h00;
    ff_ram[12615] = 8'h00;
    ff_ram[12616] = 8'h00;
    ff_ram[12617] = 8'h00;
    ff_ram[12618] = 8'h00;
    ff_ram[12619] = 8'h00;
    ff_ram[12620] = 8'h00;
    ff_ram[12621] = 8'h00;
    ff_ram[12622] = 8'h00;
    ff_ram[12623] = 8'h00;
    ff_ram[12624] = 8'h00;
    ff_ram[12625] = 8'h00;
    ff_ram[12626] = 8'h00;
    ff_ram[12627] = 8'h00;
    ff_ram[12628] = 8'h00;
    ff_ram[12629] = 8'h00;
    ff_ram[12630] = 8'h00;
    ff_ram[12631] = 8'h00;
    ff_ram[12632] = 8'h00;
    ff_ram[12633] = 8'h00;
    ff_ram[12634] = 8'h00;
    ff_ram[12635] = 8'h00;
    ff_ram[12636] = 8'h00;
    ff_ram[12637] = 8'h00;
    ff_ram[12638] = 8'h00;
    ff_ram[12639] = 8'h00;
    ff_ram[12640] = 8'h00;
    ff_ram[12641] = 8'h00;
    ff_ram[12642] = 8'h00;
    ff_ram[12643] = 8'h00;
    ff_ram[12644] = 8'h00;
    ff_ram[12645] = 8'h00;
    ff_ram[12646] = 8'h00;
    ff_ram[12647] = 8'h00;
    ff_ram[12648] = 8'h00;
    ff_ram[12649] = 8'h00;
    ff_ram[12650] = 8'h00;
    ff_ram[12651] = 8'h00;
    ff_ram[12652] = 8'h00;
    ff_ram[12653] = 8'h00;
    ff_ram[12654] = 8'h00;
    ff_ram[12655] = 8'h00;
    ff_ram[12656] = 8'h00;
    ff_ram[12657] = 8'h00;
    ff_ram[12658] = 8'h00;
    ff_ram[12659] = 8'h00;
    ff_ram[12660] = 8'h00;
    ff_ram[12661] = 8'h00;
    ff_ram[12662] = 8'h00;
    ff_ram[12663] = 8'h00;
    ff_ram[12664] = 8'h00;
    ff_ram[12665] = 8'h00;
    ff_ram[12666] = 8'h00;
    ff_ram[12667] = 8'h00;
    ff_ram[12668] = 8'h00;
    ff_ram[12669] = 8'h00;
    ff_ram[12670] = 8'h00;
    ff_ram[12671] = 8'h00;
    ff_ram[12672] = 8'h00;
    ff_ram[12673] = 8'h00;
    ff_ram[12674] = 8'h00;
    ff_ram[12675] = 8'h00;
    ff_ram[12676] = 8'h00;
    ff_ram[12677] = 8'h00;
    ff_ram[12678] = 8'h00;
    ff_ram[12679] = 8'h00;
    ff_ram[12680] = 8'h00;
    ff_ram[12681] = 8'h00;
    ff_ram[12682] = 8'h00;
    ff_ram[12683] = 8'h00;
    ff_ram[12684] = 8'h00;
    ff_ram[12685] = 8'h00;
    ff_ram[12686] = 8'h00;
    ff_ram[12687] = 8'h00;
    ff_ram[12688] = 8'h00;
    ff_ram[12689] = 8'h00;
    ff_ram[12690] = 8'h00;
    ff_ram[12691] = 8'h00;
    ff_ram[12692] = 8'h00;
    ff_ram[12693] = 8'h00;
    ff_ram[12694] = 8'h00;
    ff_ram[12695] = 8'h00;
    ff_ram[12696] = 8'h00;
    ff_ram[12697] = 8'h00;
    ff_ram[12698] = 8'h00;
    ff_ram[12699] = 8'h00;
    ff_ram[12700] = 8'h00;
    ff_ram[12701] = 8'h00;
    ff_ram[12702] = 8'h00;
    ff_ram[12703] = 8'h00;
    ff_ram[12704] = 8'h00;
    ff_ram[12705] = 8'h00;
    ff_ram[12706] = 8'h00;
    ff_ram[12707] = 8'h00;
    ff_ram[12708] = 8'h00;
    ff_ram[12709] = 8'h00;
    ff_ram[12710] = 8'h00;
    ff_ram[12711] = 8'h00;
    ff_ram[12712] = 8'h00;
    ff_ram[12713] = 8'h00;
    ff_ram[12714] = 8'h00;
    ff_ram[12715] = 8'h00;
    ff_ram[12716] = 8'h00;
    ff_ram[12717] = 8'h00;
    ff_ram[12718] = 8'h00;
    ff_ram[12719] = 8'h00;
    ff_ram[12720] = 8'h00;
    ff_ram[12721] = 8'h00;
    ff_ram[12722] = 8'h00;
    ff_ram[12723] = 8'h00;
    ff_ram[12724] = 8'h00;
    ff_ram[12725] = 8'h00;
    ff_ram[12726] = 8'h00;
    ff_ram[12727] = 8'h00;
    ff_ram[12728] = 8'h00;
    ff_ram[12729] = 8'h00;
    ff_ram[12730] = 8'h00;
    ff_ram[12731] = 8'h00;
    ff_ram[12732] = 8'h00;
    ff_ram[12733] = 8'h00;
    ff_ram[12734] = 8'h00;
    ff_ram[12735] = 8'h00;
    ff_ram[12736] = 8'h00;
    ff_ram[12737] = 8'h00;
    ff_ram[12738] = 8'h00;
    ff_ram[12739] = 8'h00;
    ff_ram[12740] = 8'h00;
    ff_ram[12741] = 8'h00;
    ff_ram[12742] = 8'h00;
    ff_ram[12743] = 8'h00;
    ff_ram[12744] = 8'h00;
    ff_ram[12745] = 8'h00;
    ff_ram[12746] = 8'h00;
    ff_ram[12747] = 8'h00;
    ff_ram[12748] = 8'h00;
    ff_ram[12749] = 8'h00;
    ff_ram[12750] = 8'h00;
    ff_ram[12751] = 8'h00;
    ff_ram[12752] = 8'h00;
    ff_ram[12753] = 8'h00;
    ff_ram[12754] = 8'h00;
    ff_ram[12755] = 8'h00;
    ff_ram[12756] = 8'h00;
    ff_ram[12757] = 8'h00;
    ff_ram[12758] = 8'h00;
    ff_ram[12759] = 8'h00;
    ff_ram[12760] = 8'h00;
    ff_ram[12761] = 8'h00;
    ff_ram[12762] = 8'h00;
    ff_ram[12763] = 8'h00;
    ff_ram[12764] = 8'h00;
    ff_ram[12765] = 8'h00;
    ff_ram[12766] = 8'h00;
    ff_ram[12767] = 8'h00;
    ff_ram[12768] = 8'h00;
    ff_ram[12769] = 8'h00;
    ff_ram[12770] = 8'h00;
    ff_ram[12771] = 8'h00;
    ff_ram[12772] = 8'h00;
    ff_ram[12773] = 8'h00;
    ff_ram[12774] = 8'h00;
    ff_ram[12775] = 8'h00;
    ff_ram[12776] = 8'h00;
    ff_ram[12777] = 8'h00;
    ff_ram[12778] = 8'h00;
    ff_ram[12779] = 8'h00;
    ff_ram[12780] = 8'h00;
    ff_ram[12781] = 8'h00;
    ff_ram[12782] = 8'h00;
    ff_ram[12783] = 8'h00;
    ff_ram[12784] = 8'h00;
    ff_ram[12785] = 8'h00;
    ff_ram[12786] = 8'h00;
    ff_ram[12787] = 8'h00;
    ff_ram[12788] = 8'h00;
    ff_ram[12789] = 8'h00;
    ff_ram[12790] = 8'h00;
    ff_ram[12791] = 8'h00;
    ff_ram[12792] = 8'h00;
    ff_ram[12793] = 8'h00;
    ff_ram[12794] = 8'h00;
    ff_ram[12795] = 8'h00;
    ff_ram[12796] = 8'h00;
    ff_ram[12797] = 8'h00;
    ff_ram[12798] = 8'h00;
    ff_ram[12799] = 8'h00;
    ff_ram[12800] = 8'h00;
    ff_ram[12801] = 8'h00;
    ff_ram[12802] = 8'h00;
    ff_ram[12803] = 8'h00;
    ff_ram[12804] = 8'h00;
    ff_ram[12805] = 8'h00;
    ff_ram[12806] = 8'h00;
    ff_ram[12807] = 8'h00;
    ff_ram[12808] = 8'h00;
    ff_ram[12809] = 8'h00;
    ff_ram[12810] = 8'h00;
    ff_ram[12811] = 8'h00;
    ff_ram[12812] = 8'h00;
    ff_ram[12813] = 8'h00;
    ff_ram[12814] = 8'h00;
    ff_ram[12815] = 8'h00;
    ff_ram[12816] = 8'h00;
    ff_ram[12817] = 8'h00;
    ff_ram[12818] = 8'h00;
    ff_ram[12819] = 8'h00;
    ff_ram[12820] = 8'h00;
    ff_ram[12821] = 8'h00;
    ff_ram[12822] = 8'h00;
    ff_ram[12823] = 8'h00;
    ff_ram[12824] = 8'h00;
    ff_ram[12825] = 8'h00;
    ff_ram[12826] = 8'h00;
    ff_ram[12827] = 8'h00;
    ff_ram[12828] = 8'h00;
    ff_ram[12829] = 8'h00;
    ff_ram[12830] = 8'h00;
    ff_ram[12831] = 8'h00;
    ff_ram[12832] = 8'h00;
    ff_ram[12833] = 8'h00;
    ff_ram[12834] = 8'h00;
    ff_ram[12835] = 8'h00;
    ff_ram[12836] = 8'h00;
    ff_ram[12837] = 8'h00;
    ff_ram[12838] = 8'h00;
    ff_ram[12839] = 8'h00;
    ff_ram[12840] = 8'h00;
    ff_ram[12841] = 8'h00;
    ff_ram[12842] = 8'h00;
    ff_ram[12843] = 8'h00;
    ff_ram[12844] = 8'h00;
    ff_ram[12845] = 8'h00;
    ff_ram[12846] = 8'h00;
    ff_ram[12847] = 8'h00;
    ff_ram[12848] = 8'h00;
    ff_ram[12849] = 8'h00;
    ff_ram[12850] = 8'h00;
    ff_ram[12851] = 8'h00;
    ff_ram[12852] = 8'h00;
    ff_ram[12853] = 8'h00;
    ff_ram[12854] = 8'h00;
    ff_ram[12855] = 8'h00;
    ff_ram[12856] = 8'h00;
    ff_ram[12857] = 8'h00;
    ff_ram[12858] = 8'h00;
    ff_ram[12859] = 8'h00;
    ff_ram[12860] = 8'h00;
    ff_ram[12861] = 8'h00;
    ff_ram[12862] = 8'h00;
    ff_ram[12863] = 8'h00;
    ff_ram[12864] = 8'h00;
    ff_ram[12865] = 8'h00;
    ff_ram[12866] = 8'h00;
    ff_ram[12867] = 8'h00;
    ff_ram[12868] = 8'h00;
    ff_ram[12869] = 8'h00;
    ff_ram[12870] = 8'h00;
    ff_ram[12871] = 8'h00;
    ff_ram[12872] = 8'h00;
    ff_ram[12873] = 8'h00;
    ff_ram[12874] = 8'h00;
    ff_ram[12875] = 8'h00;
    ff_ram[12876] = 8'h00;
    ff_ram[12877] = 8'h00;
    ff_ram[12878] = 8'h00;
    ff_ram[12879] = 8'h00;
    ff_ram[12880] = 8'h00;
    ff_ram[12881] = 8'h00;
    ff_ram[12882] = 8'h00;
    ff_ram[12883] = 8'h00;
    ff_ram[12884] = 8'h00;
    ff_ram[12885] = 8'h00;
    ff_ram[12886] = 8'h00;
    ff_ram[12887] = 8'h00;
    ff_ram[12888] = 8'h00;
    ff_ram[12889] = 8'h00;
    ff_ram[12890] = 8'h00;
    ff_ram[12891] = 8'h00;
    ff_ram[12892] = 8'h00;
    ff_ram[12893] = 8'h00;
    ff_ram[12894] = 8'h00;
    ff_ram[12895] = 8'h00;
    ff_ram[12896] = 8'h00;
    ff_ram[12897] = 8'h00;
    ff_ram[12898] = 8'h00;
    ff_ram[12899] = 8'h00;
    ff_ram[12900] = 8'h00;
    ff_ram[12901] = 8'h00;
    ff_ram[12902] = 8'h00;
    ff_ram[12903] = 8'h00;
    ff_ram[12904] = 8'h00;
    ff_ram[12905] = 8'h00;
    ff_ram[12906] = 8'h00;
    ff_ram[12907] = 8'h00;
    ff_ram[12908] = 8'h00;
    ff_ram[12909] = 8'h00;
    ff_ram[12910] = 8'h00;
    ff_ram[12911] = 8'h00;
    ff_ram[12912] = 8'h00;
    ff_ram[12913] = 8'h00;
    ff_ram[12914] = 8'h00;
    ff_ram[12915] = 8'h00;
    ff_ram[12916] = 8'h00;
    ff_ram[12917] = 8'h00;
    ff_ram[12918] = 8'h00;
    ff_ram[12919] = 8'h00;
    ff_ram[12920] = 8'h00;
    ff_ram[12921] = 8'h00;
    ff_ram[12922] = 8'h00;
    ff_ram[12923] = 8'h00;
    ff_ram[12924] = 8'h00;
    ff_ram[12925] = 8'h00;
    ff_ram[12926] = 8'h00;
    ff_ram[12927] = 8'h00;
    ff_ram[12928] = 8'h00;
    ff_ram[12929] = 8'h00;
    ff_ram[12930] = 8'h00;
    ff_ram[12931] = 8'h00;
    ff_ram[12932] = 8'h00;
    ff_ram[12933] = 8'h00;
    ff_ram[12934] = 8'h00;
    ff_ram[12935] = 8'h00;
    ff_ram[12936] = 8'h00;
    ff_ram[12937] = 8'h00;
    ff_ram[12938] = 8'h00;
    ff_ram[12939] = 8'h00;
    ff_ram[12940] = 8'h00;
    ff_ram[12941] = 8'h00;
    ff_ram[12942] = 8'h00;
    ff_ram[12943] = 8'h00;
    ff_ram[12944] = 8'h00;
    ff_ram[12945] = 8'h00;
    ff_ram[12946] = 8'h00;
    ff_ram[12947] = 8'h00;
    ff_ram[12948] = 8'h00;
    ff_ram[12949] = 8'h00;
    ff_ram[12950] = 8'h00;
    ff_ram[12951] = 8'h00;
    ff_ram[12952] = 8'h00;
    ff_ram[12953] = 8'h00;
    ff_ram[12954] = 8'h00;
    ff_ram[12955] = 8'h00;
    ff_ram[12956] = 8'h00;
    ff_ram[12957] = 8'h00;
    ff_ram[12958] = 8'h00;
    ff_ram[12959] = 8'h00;
    ff_ram[12960] = 8'h00;
    ff_ram[12961] = 8'h00;
    ff_ram[12962] = 8'h00;
    ff_ram[12963] = 8'h00;
    ff_ram[12964] = 8'h00;
    ff_ram[12965] = 8'h00;
    ff_ram[12966] = 8'h00;
    ff_ram[12967] = 8'h00;
    ff_ram[12968] = 8'h00;
    ff_ram[12969] = 8'h00;
    ff_ram[12970] = 8'h00;
    ff_ram[12971] = 8'h00;
    ff_ram[12972] = 8'h00;
    ff_ram[12973] = 8'h00;
    ff_ram[12974] = 8'h00;
    ff_ram[12975] = 8'h00;
    ff_ram[12976] = 8'h00;
    ff_ram[12977] = 8'h00;
    ff_ram[12978] = 8'h00;
    ff_ram[12979] = 8'h00;
    ff_ram[12980] = 8'h00;
    ff_ram[12981] = 8'h00;
    ff_ram[12982] = 8'h00;
    ff_ram[12983] = 8'h00;
    ff_ram[12984] = 8'h00;
    ff_ram[12985] = 8'h00;
    ff_ram[12986] = 8'h00;
    ff_ram[12987] = 8'h00;
    ff_ram[12988] = 8'h00;
    ff_ram[12989] = 8'h00;
    ff_ram[12990] = 8'h00;
    ff_ram[12991] = 8'h00;
    ff_ram[12992] = 8'h00;
    ff_ram[12993] = 8'h00;
    ff_ram[12994] = 8'h00;
    ff_ram[12995] = 8'h00;
    ff_ram[12996] = 8'h00;
    ff_ram[12997] = 8'h00;
    ff_ram[12998] = 8'h00;
    ff_ram[12999] = 8'h00;
    ff_ram[13000] = 8'h00;
    ff_ram[13001] = 8'h00;
    ff_ram[13002] = 8'h00;
    ff_ram[13003] = 8'h00;
    ff_ram[13004] = 8'h00;
    ff_ram[13005] = 8'h00;
    ff_ram[13006] = 8'h00;
    ff_ram[13007] = 8'h00;
    ff_ram[13008] = 8'h00;
    ff_ram[13009] = 8'h00;
    ff_ram[13010] = 8'h00;
    ff_ram[13011] = 8'h00;
    ff_ram[13012] = 8'h00;
    ff_ram[13013] = 8'h00;
    ff_ram[13014] = 8'h00;
    ff_ram[13015] = 8'h00;
    ff_ram[13016] = 8'h00;
    ff_ram[13017] = 8'h00;
    ff_ram[13018] = 8'h00;
    ff_ram[13019] = 8'h00;
    ff_ram[13020] = 8'h00;
    ff_ram[13021] = 8'h00;
    ff_ram[13022] = 8'h00;
    ff_ram[13023] = 8'h00;
    ff_ram[13024] = 8'h00;
    ff_ram[13025] = 8'h00;
    ff_ram[13026] = 8'h00;
    ff_ram[13027] = 8'h00;
    ff_ram[13028] = 8'h00;
    ff_ram[13029] = 8'h00;
    ff_ram[13030] = 8'h00;
    ff_ram[13031] = 8'h00;
    ff_ram[13032] = 8'h00;
    ff_ram[13033] = 8'h00;
    ff_ram[13034] = 8'h00;
    ff_ram[13035] = 8'h00;
    ff_ram[13036] = 8'h00;
    ff_ram[13037] = 8'h00;
    ff_ram[13038] = 8'h00;
    ff_ram[13039] = 8'h00;
    ff_ram[13040] = 8'h00;
    ff_ram[13041] = 8'h00;
    ff_ram[13042] = 8'h00;
    ff_ram[13043] = 8'h00;
    ff_ram[13044] = 8'h00;
    ff_ram[13045] = 8'h00;
    ff_ram[13046] = 8'h00;
    ff_ram[13047] = 8'h00;
    ff_ram[13048] = 8'h00;
    ff_ram[13049] = 8'h00;
    ff_ram[13050] = 8'h00;
    ff_ram[13051] = 8'h00;
    ff_ram[13052] = 8'h00;
    ff_ram[13053] = 8'h00;
    ff_ram[13054] = 8'h00;
    ff_ram[13055] = 8'h00;
    ff_ram[13056] = 8'h00;
    ff_ram[13057] = 8'h00;
    ff_ram[13058] = 8'h00;
    ff_ram[13059] = 8'h00;
    ff_ram[13060] = 8'h00;
    ff_ram[13061] = 8'h00;
    ff_ram[13062] = 8'h00;
    ff_ram[13063] = 8'h00;
    ff_ram[13064] = 8'h00;
    ff_ram[13065] = 8'h00;
    ff_ram[13066] = 8'h00;
    ff_ram[13067] = 8'h00;
    ff_ram[13068] = 8'h00;
    ff_ram[13069] = 8'h00;
    ff_ram[13070] = 8'h00;
    ff_ram[13071] = 8'h00;
    ff_ram[13072] = 8'h00;
    ff_ram[13073] = 8'h00;
    ff_ram[13074] = 8'h00;
    ff_ram[13075] = 8'h00;
    ff_ram[13076] = 8'h00;
    ff_ram[13077] = 8'h00;
    ff_ram[13078] = 8'h00;
    ff_ram[13079] = 8'h00;
    ff_ram[13080] = 8'h00;
    ff_ram[13081] = 8'h00;
    ff_ram[13082] = 8'h00;
    ff_ram[13083] = 8'h00;
    ff_ram[13084] = 8'h00;
    ff_ram[13085] = 8'h00;
    ff_ram[13086] = 8'h00;
    ff_ram[13087] = 8'h00;
    ff_ram[13088] = 8'h00;
    ff_ram[13089] = 8'h00;
    ff_ram[13090] = 8'h00;
    ff_ram[13091] = 8'h00;
    ff_ram[13092] = 8'h00;
    ff_ram[13093] = 8'h00;
    ff_ram[13094] = 8'h00;
    ff_ram[13095] = 8'h00;
    ff_ram[13096] = 8'h00;
    ff_ram[13097] = 8'h00;
    ff_ram[13098] = 8'h00;
    ff_ram[13099] = 8'h00;
    ff_ram[13100] = 8'h00;
    ff_ram[13101] = 8'h00;
    ff_ram[13102] = 8'h00;
    ff_ram[13103] = 8'h00;
    ff_ram[13104] = 8'h00;
    ff_ram[13105] = 8'h00;
    ff_ram[13106] = 8'h00;
    ff_ram[13107] = 8'h00;
    ff_ram[13108] = 8'h00;
    ff_ram[13109] = 8'h00;
    ff_ram[13110] = 8'h00;
    ff_ram[13111] = 8'h00;
    ff_ram[13112] = 8'h00;
    ff_ram[13113] = 8'h00;
    ff_ram[13114] = 8'h00;
    ff_ram[13115] = 8'h00;
    ff_ram[13116] = 8'h00;
    ff_ram[13117] = 8'h00;
    ff_ram[13118] = 8'h00;
    ff_ram[13119] = 8'h00;
    ff_ram[13120] = 8'h00;
    ff_ram[13121] = 8'h00;
    ff_ram[13122] = 8'h00;
    ff_ram[13123] = 8'h00;
    ff_ram[13124] = 8'h00;
    ff_ram[13125] = 8'h00;
    ff_ram[13126] = 8'h00;
    ff_ram[13127] = 8'h00;
    ff_ram[13128] = 8'h00;
    ff_ram[13129] = 8'h00;
    ff_ram[13130] = 8'h00;
    ff_ram[13131] = 8'h00;
    ff_ram[13132] = 8'h00;
    ff_ram[13133] = 8'h00;
    ff_ram[13134] = 8'h00;
    ff_ram[13135] = 8'h00;
    ff_ram[13136] = 8'h00;
    ff_ram[13137] = 8'h00;
    ff_ram[13138] = 8'h00;
    ff_ram[13139] = 8'h00;
    ff_ram[13140] = 8'h00;
    ff_ram[13141] = 8'h00;
    ff_ram[13142] = 8'h00;
    ff_ram[13143] = 8'h00;
    ff_ram[13144] = 8'h00;
    ff_ram[13145] = 8'h00;
    ff_ram[13146] = 8'h00;
    ff_ram[13147] = 8'h00;
    ff_ram[13148] = 8'h00;
    ff_ram[13149] = 8'h00;
    ff_ram[13150] = 8'h00;
    ff_ram[13151] = 8'h00;
    ff_ram[13152] = 8'h00;
    ff_ram[13153] = 8'h00;
    ff_ram[13154] = 8'h00;
    ff_ram[13155] = 8'h00;
    ff_ram[13156] = 8'h00;
    ff_ram[13157] = 8'h00;
    ff_ram[13158] = 8'h00;
    ff_ram[13159] = 8'h00;
    ff_ram[13160] = 8'h00;
    ff_ram[13161] = 8'h00;
    ff_ram[13162] = 8'h00;
    ff_ram[13163] = 8'h00;
    ff_ram[13164] = 8'h00;
    ff_ram[13165] = 8'h00;
    ff_ram[13166] = 8'h00;
    ff_ram[13167] = 8'h00;
    ff_ram[13168] = 8'h00;
    ff_ram[13169] = 8'h00;
    ff_ram[13170] = 8'h00;
    ff_ram[13171] = 8'h00;
    ff_ram[13172] = 8'h00;
    ff_ram[13173] = 8'h00;
    ff_ram[13174] = 8'h00;
    ff_ram[13175] = 8'h00;
    ff_ram[13176] = 8'h00;
    ff_ram[13177] = 8'h00;
    ff_ram[13178] = 8'h00;
    ff_ram[13179] = 8'h00;
    ff_ram[13180] = 8'h00;
    ff_ram[13181] = 8'h00;
    ff_ram[13182] = 8'h00;
    ff_ram[13183] = 8'h00;
    ff_ram[13184] = 8'h00;
    ff_ram[13185] = 8'h00;
    ff_ram[13186] = 8'h00;
    ff_ram[13187] = 8'h00;
    ff_ram[13188] = 8'h00;
    ff_ram[13189] = 8'h00;
    ff_ram[13190] = 8'h00;
    ff_ram[13191] = 8'h00;
    ff_ram[13192] = 8'h00;
    ff_ram[13193] = 8'h00;
    ff_ram[13194] = 8'h00;
    ff_ram[13195] = 8'h00;
    ff_ram[13196] = 8'h00;
    ff_ram[13197] = 8'h00;
    ff_ram[13198] = 8'h00;
    ff_ram[13199] = 8'h00;
    ff_ram[13200] = 8'h00;
    ff_ram[13201] = 8'h00;
    ff_ram[13202] = 8'h00;
    ff_ram[13203] = 8'h00;
    ff_ram[13204] = 8'h00;
    ff_ram[13205] = 8'h00;
    ff_ram[13206] = 8'h00;
    ff_ram[13207] = 8'h00;
    ff_ram[13208] = 8'h00;
    ff_ram[13209] = 8'h00;
    ff_ram[13210] = 8'h00;
    ff_ram[13211] = 8'h00;
    ff_ram[13212] = 8'h00;
    ff_ram[13213] = 8'h00;
    ff_ram[13214] = 8'h00;
    ff_ram[13215] = 8'h00;
    ff_ram[13216] = 8'h00;
    ff_ram[13217] = 8'h00;
    ff_ram[13218] = 8'h00;
    ff_ram[13219] = 8'h00;
    ff_ram[13220] = 8'h00;
    ff_ram[13221] = 8'h00;
    ff_ram[13222] = 8'h00;
    ff_ram[13223] = 8'h00;
    ff_ram[13224] = 8'h00;
    ff_ram[13225] = 8'h00;
    ff_ram[13226] = 8'h00;
    ff_ram[13227] = 8'h00;
    ff_ram[13228] = 8'h00;
    ff_ram[13229] = 8'h00;
    ff_ram[13230] = 8'h00;
    ff_ram[13231] = 8'h00;
    ff_ram[13232] = 8'h00;
    ff_ram[13233] = 8'h00;
    ff_ram[13234] = 8'h00;
    ff_ram[13235] = 8'h00;
    ff_ram[13236] = 8'h00;
    ff_ram[13237] = 8'h00;
    ff_ram[13238] = 8'h00;
    ff_ram[13239] = 8'h00;
    ff_ram[13240] = 8'h00;
    ff_ram[13241] = 8'h00;
    ff_ram[13242] = 8'h00;
    ff_ram[13243] = 8'h00;
    ff_ram[13244] = 8'h00;
    ff_ram[13245] = 8'h00;
    ff_ram[13246] = 8'h00;
    ff_ram[13247] = 8'h00;
    ff_ram[13248] = 8'h00;
    ff_ram[13249] = 8'h00;
    ff_ram[13250] = 8'h00;
    ff_ram[13251] = 8'h00;
    ff_ram[13252] = 8'h00;
    ff_ram[13253] = 8'h00;
    ff_ram[13254] = 8'h00;
    ff_ram[13255] = 8'h00;
    ff_ram[13256] = 8'h00;
    ff_ram[13257] = 8'h00;
    ff_ram[13258] = 8'h00;
    ff_ram[13259] = 8'h00;
    ff_ram[13260] = 8'h00;
    ff_ram[13261] = 8'h00;
    ff_ram[13262] = 8'h00;
    ff_ram[13263] = 8'h00;
    ff_ram[13264] = 8'h00;
    ff_ram[13265] = 8'h00;
    ff_ram[13266] = 8'h00;
    ff_ram[13267] = 8'h00;
    ff_ram[13268] = 8'h00;
    ff_ram[13269] = 8'h00;
    ff_ram[13270] = 8'h00;
    ff_ram[13271] = 8'h00;
    ff_ram[13272] = 8'h00;
    ff_ram[13273] = 8'h00;
    ff_ram[13274] = 8'h00;
    ff_ram[13275] = 8'h00;
    ff_ram[13276] = 8'h00;
    ff_ram[13277] = 8'h00;
    ff_ram[13278] = 8'h00;
    ff_ram[13279] = 8'h00;
    ff_ram[13280] = 8'h00;
    ff_ram[13281] = 8'h00;
    ff_ram[13282] = 8'h00;
    ff_ram[13283] = 8'h00;
    ff_ram[13284] = 8'h00;
    ff_ram[13285] = 8'h00;
    ff_ram[13286] = 8'h00;
    ff_ram[13287] = 8'h00;
    ff_ram[13288] = 8'h00;
    ff_ram[13289] = 8'h00;
    ff_ram[13290] = 8'h00;
    ff_ram[13291] = 8'h00;
    ff_ram[13292] = 8'h00;
    ff_ram[13293] = 8'h00;
    ff_ram[13294] = 8'h00;
    ff_ram[13295] = 8'h00;
    ff_ram[13296] = 8'h00;
    ff_ram[13297] = 8'h00;
    ff_ram[13298] = 8'h00;
    ff_ram[13299] = 8'h00;
    ff_ram[13300] = 8'h00;
    ff_ram[13301] = 8'h00;
    ff_ram[13302] = 8'h00;
    ff_ram[13303] = 8'h00;
    ff_ram[13304] = 8'h00;
    ff_ram[13305] = 8'h00;
    ff_ram[13306] = 8'h00;
    ff_ram[13307] = 8'h00;
    ff_ram[13308] = 8'h00;
    ff_ram[13309] = 8'h00;
    ff_ram[13310] = 8'h00;
    ff_ram[13311] = 8'h00;
    ff_ram[13312] = 8'h00;
    ff_ram[13313] = 8'h00;
    ff_ram[13314] = 8'h00;
    ff_ram[13315] = 8'h00;
    ff_ram[13316] = 8'h00;
    ff_ram[13317] = 8'h00;
    ff_ram[13318] = 8'h00;
    ff_ram[13319] = 8'h00;
    ff_ram[13320] = 8'h00;
    ff_ram[13321] = 8'h00;
    ff_ram[13322] = 8'h00;
    ff_ram[13323] = 8'h00;
    ff_ram[13324] = 8'h00;
    ff_ram[13325] = 8'h00;
    ff_ram[13326] = 8'h00;
    ff_ram[13327] = 8'h00;
    ff_ram[13328] = 8'h00;
    ff_ram[13329] = 8'h00;
    ff_ram[13330] = 8'h00;
    ff_ram[13331] = 8'h00;
    ff_ram[13332] = 8'h00;
    ff_ram[13333] = 8'h00;
    ff_ram[13334] = 8'h00;
    ff_ram[13335] = 8'h00;
    ff_ram[13336] = 8'h00;
    ff_ram[13337] = 8'h00;
    ff_ram[13338] = 8'h00;
    ff_ram[13339] = 8'h00;
    ff_ram[13340] = 8'h00;
    ff_ram[13341] = 8'h00;
    ff_ram[13342] = 8'h00;
    ff_ram[13343] = 8'h00;
    ff_ram[13344] = 8'h00;
    ff_ram[13345] = 8'h00;
    ff_ram[13346] = 8'h00;
    ff_ram[13347] = 8'h00;
    ff_ram[13348] = 8'h00;
    ff_ram[13349] = 8'h00;
    ff_ram[13350] = 8'h00;
    ff_ram[13351] = 8'h00;
    ff_ram[13352] = 8'h00;
    ff_ram[13353] = 8'h00;
    ff_ram[13354] = 8'h00;
    ff_ram[13355] = 8'h00;
    ff_ram[13356] = 8'h00;
    ff_ram[13357] = 8'h00;
    ff_ram[13358] = 8'h00;
    ff_ram[13359] = 8'h00;
    ff_ram[13360] = 8'h00;
    ff_ram[13361] = 8'h00;
    ff_ram[13362] = 8'h00;
    ff_ram[13363] = 8'h00;
    ff_ram[13364] = 8'h00;
    ff_ram[13365] = 8'h00;
    ff_ram[13366] = 8'h00;
    ff_ram[13367] = 8'h00;
    ff_ram[13368] = 8'h00;
    ff_ram[13369] = 8'h00;
    ff_ram[13370] = 8'h00;
    ff_ram[13371] = 8'h00;
    ff_ram[13372] = 8'h00;
    ff_ram[13373] = 8'h00;
    ff_ram[13374] = 8'h00;
    ff_ram[13375] = 8'h00;
    ff_ram[13376] = 8'h00;
    ff_ram[13377] = 8'h00;
    ff_ram[13378] = 8'h00;
    ff_ram[13379] = 8'h00;
    ff_ram[13380] = 8'h00;
    ff_ram[13381] = 8'h00;
    ff_ram[13382] = 8'h00;
    ff_ram[13383] = 8'h00;
    ff_ram[13384] = 8'h00;
    ff_ram[13385] = 8'h00;
    ff_ram[13386] = 8'h00;
    ff_ram[13387] = 8'h00;
    ff_ram[13388] = 8'h00;
    ff_ram[13389] = 8'h00;
    ff_ram[13390] = 8'h00;
    ff_ram[13391] = 8'h00;
    ff_ram[13392] = 8'h00;
    ff_ram[13393] = 8'h00;
    ff_ram[13394] = 8'h00;
    ff_ram[13395] = 8'h00;
    ff_ram[13396] = 8'h00;
    ff_ram[13397] = 8'h00;
    ff_ram[13398] = 8'h00;
    ff_ram[13399] = 8'h00;
    ff_ram[13400] = 8'h00;
    ff_ram[13401] = 8'h00;
    ff_ram[13402] = 8'h00;
    ff_ram[13403] = 8'h00;
    ff_ram[13404] = 8'h00;
    ff_ram[13405] = 8'h00;
    ff_ram[13406] = 8'h00;
    ff_ram[13407] = 8'h00;
    ff_ram[13408] = 8'h00;
    ff_ram[13409] = 8'h00;
    ff_ram[13410] = 8'h00;
    ff_ram[13411] = 8'h00;
    ff_ram[13412] = 8'h00;
    ff_ram[13413] = 8'h00;
    ff_ram[13414] = 8'h00;
    ff_ram[13415] = 8'h00;
    ff_ram[13416] = 8'h00;
    ff_ram[13417] = 8'h00;
    ff_ram[13418] = 8'h00;
    ff_ram[13419] = 8'h00;
    ff_ram[13420] = 8'h00;
    ff_ram[13421] = 8'h00;
    ff_ram[13422] = 8'h00;
    ff_ram[13423] = 8'h00;
    ff_ram[13424] = 8'h00;
    ff_ram[13425] = 8'h00;
    ff_ram[13426] = 8'h00;
    ff_ram[13427] = 8'h00;
    ff_ram[13428] = 8'h00;
    ff_ram[13429] = 8'h00;
    ff_ram[13430] = 8'h00;
    ff_ram[13431] = 8'h00;
    ff_ram[13432] = 8'h00;
    ff_ram[13433] = 8'h00;
    ff_ram[13434] = 8'h00;
    ff_ram[13435] = 8'h00;
    ff_ram[13436] = 8'h00;
    ff_ram[13437] = 8'h00;
    ff_ram[13438] = 8'h00;
    ff_ram[13439] = 8'h00;
    ff_ram[13440] = 8'h00;
    ff_ram[13441] = 8'h00;
    ff_ram[13442] = 8'h00;
    ff_ram[13443] = 8'h00;
    ff_ram[13444] = 8'h00;
    ff_ram[13445] = 8'h00;
    ff_ram[13446] = 8'h00;
    ff_ram[13447] = 8'h00;
    ff_ram[13448] = 8'h00;
    ff_ram[13449] = 8'h00;
    ff_ram[13450] = 8'h00;
    ff_ram[13451] = 8'h00;
    ff_ram[13452] = 8'h00;
    ff_ram[13453] = 8'h00;
    ff_ram[13454] = 8'h00;
    ff_ram[13455] = 8'h00;
    ff_ram[13456] = 8'h00;
    ff_ram[13457] = 8'h00;
    ff_ram[13458] = 8'h00;
    ff_ram[13459] = 8'h00;
    ff_ram[13460] = 8'h00;
    ff_ram[13461] = 8'h00;
    ff_ram[13462] = 8'h00;
    ff_ram[13463] = 8'h00;
    ff_ram[13464] = 8'h00;
    ff_ram[13465] = 8'h00;
    ff_ram[13466] = 8'h00;
    ff_ram[13467] = 8'h00;
    ff_ram[13468] = 8'h00;
    ff_ram[13469] = 8'h00;
    ff_ram[13470] = 8'h00;
    ff_ram[13471] = 8'h00;
    ff_ram[13472] = 8'h00;
    ff_ram[13473] = 8'h00;
    ff_ram[13474] = 8'h00;
    ff_ram[13475] = 8'h00;
    ff_ram[13476] = 8'h00;
    ff_ram[13477] = 8'h00;
    ff_ram[13478] = 8'h00;
    ff_ram[13479] = 8'h00;
    ff_ram[13480] = 8'h00;
    ff_ram[13481] = 8'h00;
    ff_ram[13482] = 8'h00;
    ff_ram[13483] = 8'h00;
    ff_ram[13484] = 8'h00;
    ff_ram[13485] = 8'h00;
    ff_ram[13486] = 8'h00;
    ff_ram[13487] = 8'h00;
    ff_ram[13488] = 8'h00;
    ff_ram[13489] = 8'h00;
    ff_ram[13490] = 8'h00;
    ff_ram[13491] = 8'h00;
    ff_ram[13492] = 8'h00;
    ff_ram[13493] = 8'h00;
    ff_ram[13494] = 8'h00;
    ff_ram[13495] = 8'h00;
    ff_ram[13496] = 8'h00;
    ff_ram[13497] = 8'h00;
    ff_ram[13498] = 8'h00;
    ff_ram[13499] = 8'h00;
    ff_ram[13500] = 8'h00;
    ff_ram[13501] = 8'h00;
    ff_ram[13502] = 8'h00;
    ff_ram[13503] = 8'h00;
    ff_ram[13504] = 8'h00;
    ff_ram[13505] = 8'h00;
    ff_ram[13506] = 8'h00;
    ff_ram[13507] = 8'h00;
    ff_ram[13508] = 8'h00;
    ff_ram[13509] = 8'h00;
    ff_ram[13510] = 8'h00;
    ff_ram[13511] = 8'h00;
    ff_ram[13512] = 8'h00;
    ff_ram[13513] = 8'h00;
    ff_ram[13514] = 8'h00;
    ff_ram[13515] = 8'h00;
    ff_ram[13516] = 8'h00;
    ff_ram[13517] = 8'h00;
    ff_ram[13518] = 8'h00;
    ff_ram[13519] = 8'h00;
    ff_ram[13520] = 8'h00;
    ff_ram[13521] = 8'h00;
    ff_ram[13522] = 8'h00;
    ff_ram[13523] = 8'h00;
    ff_ram[13524] = 8'h00;
    ff_ram[13525] = 8'h00;
    ff_ram[13526] = 8'h00;
    ff_ram[13527] = 8'h00;
    ff_ram[13528] = 8'h00;
    ff_ram[13529] = 8'h00;
    ff_ram[13530] = 8'h00;
    ff_ram[13531] = 8'h00;
    ff_ram[13532] = 8'h00;
    ff_ram[13533] = 8'h00;
    ff_ram[13534] = 8'h00;
    ff_ram[13535] = 8'h00;
    ff_ram[13536] = 8'h00;
    ff_ram[13537] = 8'h00;
    ff_ram[13538] = 8'h00;
    ff_ram[13539] = 8'h00;
    ff_ram[13540] = 8'h00;
    ff_ram[13541] = 8'h00;
    ff_ram[13542] = 8'h00;
    ff_ram[13543] = 8'h00;
    ff_ram[13544] = 8'h00;
    ff_ram[13545] = 8'h00;
    ff_ram[13546] = 8'h00;
    ff_ram[13547] = 8'h00;
    ff_ram[13548] = 8'h00;
    ff_ram[13549] = 8'h00;
    ff_ram[13550] = 8'h00;
    ff_ram[13551] = 8'h00;
    ff_ram[13552] = 8'h00;
    ff_ram[13553] = 8'h00;
    ff_ram[13554] = 8'h00;
    ff_ram[13555] = 8'h00;
    ff_ram[13556] = 8'h00;
    ff_ram[13557] = 8'h00;
    ff_ram[13558] = 8'h00;
    ff_ram[13559] = 8'h00;
    ff_ram[13560] = 8'h00;
    ff_ram[13561] = 8'h00;
    ff_ram[13562] = 8'h00;
    ff_ram[13563] = 8'h00;
    ff_ram[13564] = 8'h00;
    ff_ram[13565] = 8'h00;
    ff_ram[13566] = 8'h00;
    ff_ram[13567] = 8'h00;
    ff_ram[13568] = 8'h00;
    ff_ram[13569] = 8'h00;
    ff_ram[13570] = 8'h00;
    ff_ram[13571] = 8'h00;
    ff_ram[13572] = 8'h00;
    ff_ram[13573] = 8'h00;
    ff_ram[13574] = 8'h00;
    ff_ram[13575] = 8'h00;
    ff_ram[13576] = 8'h00;
    ff_ram[13577] = 8'h00;
    ff_ram[13578] = 8'h00;
    ff_ram[13579] = 8'h00;
    ff_ram[13580] = 8'h00;
    ff_ram[13581] = 8'h00;
    ff_ram[13582] = 8'h00;
    ff_ram[13583] = 8'h00;
    ff_ram[13584] = 8'h00;
    ff_ram[13585] = 8'h00;
    ff_ram[13586] = 8'h00;
    ff_ram[13587] = 8'h00;
    ff_ram[13588] = 8'h00;
    ff_ram[13589] = 8'h00;
    ff_ram[13590] = 8'h00;
    ff_ram[13591] = 8'h00;
    ff_ram[13592] = 8'h00;
    ff_ram[13593] = 8'h00;
    ff_ram[13594] = 8'h00;
    ff_ram[13595] = 8'h00;
    ff_ram[13596] = 8'h00;
    ff_ram[13597] = 8'h00;
    ff_ram[13598] = 8'h00;
    ff_ram[13599] = 8'h00;
    ff_ram[13600] = 8'h00;
    ff_ram[13601] = 8'h00;
    ff_ram[13602] = 8'h00;
    ff_ram[13603] = 8'h00;
    ff_ram[13604] = 8'h00;
    ff_ram[13605] = 8'h00;
    ff_ram[13606] = 8'h00;
    ff_ram[13607] = 8'h00;
    ff_ram[13608] = 8'h00;
    ff_ram[13609] = 8'h00;
    ff_ram[13610] = 8'h00;
    ff_ram[13611] = 8'h00;
    ff_ram[13612] = 8'h00;
    ff_ram[13613] = 8'h00;
    ff_ram[13614] = 8'h00;
    ff_ram[13615] = 8'h00;
    ff_ram[13616] = 8'h00;
    ff_ram[13617] = 8'h00;
    ff_ram[13618] = 8'h00;
    ff_ram[13619] = 8'h00;
    ff_ram[13620] = 8'h00;
    ff_ram[13621] = 8'h00;
    ff_ram[13622] = 8'h00;
    ff_ram[13623] = 8'h00;
    ff_ram[13624] = 8'h00;
    ff_ram[13625] = 8'h00;
    ff_ram[13626] = 8'h00;
    ff_ram[13627] = 8'h00;
    ff_ram[13628] = 8'h00;
    ff_ram[13629] = 8'h00;
    ff_ram[13630] = 8'h00;
    ff_ram[13631] = 8'h00;
    ff_ram[13632] = 8'h00;
    ff_ram[13633] = 8'h00;
    ff_ram[13634] = 8'h00;
    ff_ram[13635] = 8'h00;
    ff_ram[13636] = 8'h00;
    ff_ram[13637] = 8'h00;
    ff_ram[13638] = 8'h00;
    ff_ram[13639] = 8'h00;
    ff_ram[13640] = 8'h00;
    ff_ram[13641] = 8'h00;
    ff_ram[13642] = 8'h00;
    ff_ram[13643] = 8'h00;
    ff_ram[13644] = 8'h00;
    ff_ram[13645] = 8'h00;
    ff_ram[13646] = 8'h00;
    ff_ram[13647] = 8'h00;
    ff_ram[13648] = 8'h00;
    ff_ram[13649] = 8'h00;
    ff_ram[13650] = 8'h00;
    ff_ram[13651] = 8'h00;
    ff_ram[13652] = 8'h00;
    ff_ram[13653] = 8'h00;
    ff_ram[13654] = 8'h00;
    ff_ram[13655] = 8'h00;
    ff_ram[13656] = 8'h00;
    ff_ram[13657] = 8'h00;
    ff_ram[13658] = 8'h00;
    ff_ram[13659] = 8'h00;
    ff_ram[13660] = 8'h00;
    ff_ram[13661] = 8'h00;
    ff_ram[13662] = 8'h00;
    ff_ram[13663] = 8'h00;
    ff_ram[13664] = 8'h00;
    ff_ram[13665] = 8'h00;
    ff_ram[13666] = 8'h00;
    ff_ram[13667] = 8'h00;
    ff_ram[13668] = 8'h00;
    ff_ram[13669] = 8'h00;
    ff_ram[13670] = 8'h00;
    ff_ram[13671] = 8'h00;
    ff_ram[13672] = 8'h00;
    ff_ram[13673] = 8'h00;
    ff_ram[13674] = 8'h00;
    ff_ram[13675] = 8'h00;
    ff_ram[13676] = 8'h00;
    ff_ram[13677] = 8'h00;
    ff_ram[13678] = 8'h00;
    ff_ram[13679] = 8'h00;
    ff_ram[13680] = 8'h00;
    ff_ram[13681] = 8'h00;
    ff_ram[13682] = 8'h00;
    ff_ram[13683] = 8'h00;
    ff_ram[13684] = 8'h00;
    ff_ram[13685] = 8'h00;
    ff_ram[13686] = 8'h00;
    ff_ram[13687] = 8'h00;
    ff_ram[13688] = 8'h00;
    ff_ram[13689] = 8'h00;
    ff_ram[13690] = 8'h00;
    ff_ram[13691] = 8'h00;
    ff_ram[13692] = 8'h00;
    ff_ram[13693] = 8'h00;
    ff_ram[13694] = 8'h00;
    ff_ram[13695] = 8'h00;
    ff_ram[13696] = 8'h00;
    ff_ram[13697] = 8'h00;
    ff_ram[13698] = 8'h00;
    ff_ram[13699] = 8'h00;
    ff_ram[13700] = 8'h00;
    ff_ram[13701] = 8'h00;
    ff_ram[13702] = 8'h00;
    ff_ram[13703] = 8'h00;
    ff_ram[13704] = 8'h00;
    ff_ram[13705] = 8'h00;
    ff_ram[13706] = 8'h00;
    ff_ram[13707] = 8'h00;
    ff_ram[13708] = 8'h00;
    ff_ram[13709] = 8'h00;
    ff_ram[13710] = 8'h00;
    ff_ram[13711] = 8'h00;
    ff_ram[13712] = 8'h00;
    ff_ram[13713] = 8'h00;
    ff_ram[13714] = 8'h00;
    ff_ram[13715] = 8'h00;
    ff_ram[13716] = 8'h00;
    ff_ram[13717] = 8'h00;
    ff_ram[13718] = 8'h00;
    ff_ram[13719] = 8'h00;
    ff_ram[13720] = 8'h00;
    ff_ram[13721] = 8'h00;
    ff_ram[13722] = 8'h00;
    ff_ram[13723] = 8'h00;
    ff_ram[13724] = 8'h00;
    ff_ram[13725] = 8'h00;
    ff_ram[13726] = 8'h00;
    ff_ram[13727] = 8'h00;
    ff_ram[13728] = 8'h00;
    ff_ram[13729] = 8'h00;
    ff_ram[13730] = 8'h00;
    ff_ram[13731] = 8'h00;
    ff_ram[13732] = 8'h00;
    ff_ram[13733] = 8'h00;
    ff_ram[13734] = 8'h00;
    ff_ram[13735] = 8'h00;
    ff_ram[13736] = 8'h00;
    ff_ram[13737] = 8'h00;
    ff_ram[13738] = 8'h00;
    ff_ram[13739] = 8'h00;
    ff_ram[13740] = 8'h00;
    ff_ram[13741] = 8'h00;
    ff_ram[13742] = 8'h00;
    ff_ram[13743] = 8'h00;
    ff_ram[13744] = 8'h00;
    ff_ram[13745] = 8'h00;
    ff_ram[13746] = 8'h00;
    ff_ram[13747] = 8'h00;
    ff_ram[13748] = 8'h00;
    ff_ram[13749] = 8'h00;
    ff_ram[13750] = 8'h00;
    ff_ram[13751] = 8'h00;
    ff_ram[13752] = 8'h00;
    ff_ram[13753] = 8'h00;
    ff_ram[13754] = 8'h00;
    ff_ram[13755] = 8'h00;
    ff_ram[13756] = 8'h00;
    ff_ram[13757] = 8'h00;
    ff_ram[13758] = 8'h00;
    ff_ram[13759] = 8'h00;
    ff_ram[13760] = 8'h00;
    ff_ram[13761] = 8'h00;
    ff_ram[13762] = 8'h00;
    ff_ram[13763] = 8'h00;
    ff_ram[13764] = 8'h00;
    ff_ram[13765] = 8'h00;
    ff_ram[13766] = 8'h00;
    ff_ram[13767] = 8'h00;
    ff_ram[13768] = 8'h00;
    ff_ram[13769] = 8'h00;
    ff_ram[13770] = 8'h00;
    ff_ram[13771] = 8'h00;
    ff_ram[13772] = 8'h00;
    ff_ram[13773] = 8'h00;
    ff_ram[13774] = 8'h00;
    ff_ram[13775] = 8'h00;
    ff_ram[13776] = 8'h00;
    ff_ram[13777] = 8'h00;
    ff_ram[13778] = 8'h00;
    ff_ram[13779] = 8'h00;
    ff_ram[13780] = 8'h00;
    ff_ram[13781] = 8'h00;
    ff_ram[13782] = 8'h00;
    ff_ram[13783] = 8'h00;
    ff_ram[13784] = 8'h00;
    ff_ram[13785] = 8'h00;
    ff_ram[13786] = 8'h00;
    ff_ram[13787] = 8'h00;
    ff_ram[13788] = 8'h00;
    ff_ram[13789] = 8'h00;
    ff_ram[13790] = 8'h00;
    ff_ram[13791] = 8'h00;
    ff_ram[13792] = 8'h00;
    ff_ram[13793] = 8'h00;
    ff_ram[13794] = 8'h00;
    ff_ram[13795] = 8'h00;
    ff_ram[13796] = 8'h00;
    ff_ram[13797] = 8'h00;
    ff_ram[13798] = 8'h00;
    ff_ram[13799] = 8'h00;
    ff_ram[13800] = 8'h00;
    ff_ram[13801] = 8'h00;
    ff_ram[13802] = 8'h00;
    ff_ram[13803] = 8'h00;
    ff_ram[13804] = 8'h00;
    ff_ram[13805] = 8'h00;
    ff_ram[13806] = 8'h00;
    ff_ram[13807] = 8'h00;
    ff_ram[13808] = 8'h00;
    ff_ram[13809] = 8'h00;
    ff_ram[13810] = 8'h00;
    ff_ram[13811] = 8'h00;
    ff_ram[13812] = 8'h00;
    ff_ram[13813] = 8'h00;
    ff_ram[13814] = 8'h00;
    ff_ram[13815] = 8'h00;
    ff_ram[13816] = 8'h00;
    ff_ram[13817] = 8'h00;
    ff_ram[13818] = 8'h00;
    ff_ram[13819] = 8'h00;
    ff_ram[13820] = 8'h00;
    ff_ram[13821] = 8'h00;
    ff_ram[13822] = 8'h00;
    ff_ram[13823] = 8'h00;
    ff_ram[13824] = 8'h00;
    ff_ram[13825] = 8'h00;
    ff_ram[13826] = 8'h00;
    ff_ram[13827] = 8'h00;
    ff_ram[13828] = 8'h00;
    ff_ram[13829] = 8'h00;
    ff_ram[13830] = 8'h00;
    ff_ram[13831] = 8'h00;
    ff_ram[13832] = 8'h00;
    ff_ram[13833] = 8'h00;
    ff_ram[13834] = 8'h00;
    ff_ram[13835] = 8'h00;
    ff_ram[13836] = 8'h00;
    ff_ram[13837] = 8'h00;
    ff_ram[13838] = 8'h00;
    ff_ram[13839] = 8'h00;
    ff_ram[13840] = 8'h00;
    ff_ram[13841] = 8'h00;
    ff_ram[13842] = 8'h00;
    ff_ram[13843] = 8'h00;
    ff_ram[13844] = 8'h00;
    ff_ram[13845] = 8'h00;
    ff_ram[13846] = 8'h00;
    ff_ram[13847] = 8'h00;
    ff_ram[13848] = 8'h00;
    ff_ram[13849] = 8'h00;
    ff_ram[13850] = 8'h00;
    ff_ram[13851] = 8'h00;
    ff_ram[13852] = 8'h00;
    ff_ram[13853] = 8'h00;
    ff_ram[13854] = 8'h00;
    ff_ram[13855] = 8'h00;
    ff_ram[13856] = 8'h00;
    ff_ram[13857] = 8'h00;
    ff_ram[13858] = 8'h00;
    ff_ram[13859] = 8'h00;
    ff_ram[13860] = 8'h00;
    ff_ram[13861] = 8'h00;
    ff_ram[13862] = 8'h00;
    ff_ram[13863] = 8'h00;
    ff_ram[13864] = 8'h00;
    ff_ram[13865] = 8'h00;
    ff_ram[13866] = 8'h00;
    ff_ram[13867] = 8'h00;
    ff_ram[13868] = 8'h00;
    ff_ram[13869] = 8'h00;
    ff_ram[13870] = 8'h00;
    ff_ram[13871] = 8'h00;
    ff_ram[13872] = 8'h00;
    ff_ram[13873] = 8'h00;
    ff_ram[13874] = 8'h00;
    ff_ram[13875] = 8'h00;
    ff_ram[13876] = 8'h00;
    ff_ram[13877] = 8'h00;
    ff_ram[13878] = 8'h00;
    ff_ram[13879] = 8'h00;
    ff_ram[13880] = 8'h00;
    ff_ram[13881] = 8'h00;
    ff_ram[13882] = 8'h00;
    ff_ram[13883] = 8'h00;
    ff_ram[13884] = 8'h00;
    ff_ram[13885] = 8'h00;
    ff_ram[13886] = 8'h00;
    ff_ram[13887] = 8'h00;
    ff_ram[13888] = 8'h00;
    ff_ram[13889] = 8'h00;
    ff_ram[13890] = 8'h00;
    ff_ram[13891] = 8'h00;
    ff_ram[13892] = 8'h00;
    ff_ram[13893] = 8'h00;
    ff_ram[13894] = 8'h00;
    ff_ram[13895] = 8'h00;
    ff_ram[13896] = 8'h00;
    ff_ram[13897] = 8'h00;
    ff_ram[13898] = 8'h00;
    ff_ram[13899] = 8'h00;
    ff_ram[13900] = 8'h00;
    ff_ram[13901] = 8'h00;
    ff_ram[13902] = 8'h00;
    ff_ram[13903] = 8'h00;
    ff_ram[13904] = 8'h00;
    ff_ram[13905] = 8'h00;
    ff_ram[13906] = 8'h00;
    ff_ram[13907] = 8'h00;
    ff_ram[13908] = 8'h00;
    ff_ram[13909] = 8'h00;
    ff_ram[13910] = 8'h00;
    ff_ram[13911] = 8'h00;
    ff_ram[13912] = 8'h00;
    ff_ram[13913] = 8'h00;
    ff_ram[13914] = 8'h00;
    ff_ram[13915] = 8'h00;
    ff_ram[13916] = 8'h00;
    ff_ram[13917] = 8'h00;
    ff_ram[13918] = 8'h00;
    ff_ram[13919] = 8'h00;
    ff_ram[13920] = 8'h00;
    ff_ram[13921] = 8'h00;
    ff_ram[13922] = 8'h00;
    ff_ram[13923] = 8'h00;
    ff_ram[13924] = 8'h00;
    ff_ram[13925] = 8'h00;
    ff_ram[13926] = 8'h00;
    ff_ram[13927] = 8'h00;
    ff_ram[13928] = 8'h00;
    ff_ram[13929] = 8'h00;
    ff_ram[13930] = 8'h00;
    ff_ram[13931] = 8'h00;
    ff_ram[13932] = 8'h00;
    ff_ram[13933] = 8'h00;
    ff_ram[13934] = 8'h00;
    ff_ram[13935] = 8'h00;
    ff_ram[13936] = 8'h00;
    ff_ram[13937] = 8'h00;
    ff_ram[13938] = 8'h00;
    ff_ram[13939] = 8'h00;
    ff_ram[13940] = 8'h00;
    ff_ram[13941] = 8'h00;
    ff_ram[13942] = 8'h00;
    ff_ram[13943] = 8'h00;
    ff_ram[13944] = 8'h00;
    ff_ram[13945] = 8'h00;
    ff_ram[13946] = 8'h00;
    ff_ram[13947] = 8'h00;
    ff_ram[13948] = 8'h00;
    ff_ram[13949] = 8'h00;
    ff_ram[13950] = 8'h00;
    ff_ram[13951] = 8'h00;
    ff_ram[13952] = 8'h00;
    ff_ram[13953] = 8'h00;
    ff_ram[13954] = 8'h00;
    ff_ram[13955] = 8'h00;
    ff_ram[13956] = 8'h00;
    ff_ram[13957] = 8'h00;
    ff_ram[13958] = 8'h00;
    ff_ram[13959] = 8'h00;
    ff_ram[13960] = 8'h00;
    ff_ram[13961] = 8'h00;
    ff_ram[13962] = 8'h00;
    ff_ram[13963] = 8'h00;
    ff_ram[13964] = 8'h00;
    ff_ram[13965] = 8'h00;
    ff_ram[13966] = 8'h00;
    ff_ram[13967] = 8'h00;
    ff_ram[13968] = 8'h00;
    ff_ram[13969] = 8'h00;
    ff_ram[13970] = 8'h00;
    ff_ram[13971] = 8'h00;
    ff_ram[13972] = 8'h00;
    ff_ram[13973] = 8'h00;
    ff_ram[13974] = 8'h00;
    ff_ram[13975] = 8'h00;
    ff_ram[13976] = 8'h00;
    ff_ram[13977] = 8'h00;
    ff_ram[13978] = 8'h00;
    ff_ram[13979] = 8'h00;
    ff_ram[13980] = 8'h00;
    ff_ram[13981] = 8'h00;
    ff_ram[13982] = 8'h00;
    ff_ram[13983] = 8'h00;
    ff_ram[13984] = 8'h00;
    ff_ram[13985] = 8'h00;
    ff_ram[13986] = 8'h00;
    ff_ram[13987] = 8'h00;
    ff_ram[13988] = 8'h00;
    ff_ram[13989] = 8'h00;
    ff_ram[13990] = 8'h00;
    ff_ram[13991] = 8'h00;
    ff_ram[13992] = 8'h00;
    ff_ram[13993] = 8'h00;
    ff_ram[13994] = 8'h00;
    ff_ram[13995] = 8'h00;
    ff_ram[13996] = 8'h00;
    ff_ram[13997] = 8'h00;
    ff_ram[13998] = 8'h00;
    ff_ram[13999] = 8'h00;
    ff_ram[14000] = 8'h00;
    ff_ram[14001] = 8'h00;
    ff_ram[14002] = 8'h00;
    ff_ram[14003] = 8'h00;
    ff_ram[14004] = 8'h00;
    ff_ram[14005] = 8'h00;
    ff_ram[14006] = 8'h00;
    ff_ram[14007] = 8'h00;
    ff_ram[14008] = 8'h00;
    ff_ram[14009] = 8'h00;
    ff_ram[14010] = 8'h00;
    ff_ram[14011] = 8'h00;
    ff_ram[14012] = 8'h00;
    ff_ram[14013] = 8'h00;
    ff_ram[14014] = 8'h00;
    ff_ram[14015] = 8'h00;
    ff_ram[14016] = 8'h00;
    ff_ram[14017] = 8'h00;
    ff_ram[14018] = 8'h00;
    ff_ram[14019] = 8'h00;
    ff_ram[14020] = 8'h00;
    ff_ram[14021] = 8'h00;
    ff_ram[14022] = 8'h00;
    ff_ram[14023] = 8'h00;
    ff_ram[14024] = 8'h00;
    ff_ram[14025] = 8'h00;
    ff_ram[14026] = 8'h00;
    ff_ram[14027] = 8'h00;
    ff_ram[14028] = 8'h00;
    ff_ram[14029] = 8'h00;
    ff_ram[14030] = 8'h00;
    ff_ram[14031] = 8'h00;
    ff_ram[14032] = 8'h00;
    ff_ram[14033] = 8'h00;
    ff_ram[14034] = 8'h00;
    ff_ram[14035] = 8'h00;
    ff_ram[14036] = 8'h00;
    ff_ram[14037] = 8'h00;
    ff_ram[14038] = 8'h00;
    ff_ram[14039] = 8'h00;
    ff_ram[14040] = 8'h00;
    ff_ram[14041] = 8'h00;
    ff_ram[14042] = 8'h00;
    ff_ram[14043] = 8'h00;
    ff_ram[14044] = 8'h00;
    ff_ram[14045] = 8'h00;
    ff_ram[14046] = 8'h00;
    ff_ram[14047] = 8'h00;
    ff_ram[14048] = 8'h00;
    ff_ram[14049] = 8'h00;
    ff_ram[14050] = 8'h00;
    ff_ram[14051] = 8'h00;
    ff_ram[14052] = 8'h00;
    ff_ram[14053] = 8'h00;
    ff_ram[14054] = 8'h00;
    ff_ram[14055] = 8'h00;
    ff_ram[14056] = 8'h00;
    ff_ram[14057] = 8'h00;
    ff_ram[14058] = 8'h00;
    ff_ram[14059] = 8'h00;
    ff_ram[14060] = 8'h00;
    ff_ram[14061] = 8'h00;
    ff_ram[14062] = 8'h00;
    ff_ram[14063] = 8'h00;
    ff_ram[14064] = 8'h00;
    ff_ram[14065] = 8'h00;
    ff_ram[14066] = 8'h00;
    ff_ram[14067] = 8'h00;
    ff_ram[14068] = 8'h00;
    ff_ram[14069] = 8'h00;
    ff_ram[14070] = 8'h00;
    ff_ram[14071] = 8'h00;
    ff_ram[14072] = 8'h00;
    ff_ram[14073] = 8'h00;
    ff_ram[14074] = 8'h00;
    ff_ram[14075] = 8'h00;
    ff_ram[14076] = 8'h00;
    ff_ram[14077] = 8'h00;
    ff_ram[14078] = 8'h00;
    ff_ram[14079] = 8'h00;
    ff_ram[14080] = 8'h00;
    ff_ram[14081] = 8'h00;
    ff_ram[14082] = 8'h00;
    ff_ram[14083] = 8'h00;
    ff_ram[14084] = 8'h00;
    ff_ram[14085] = 8'h00;
    ff_ram[14086] = 8'h00;
    ff_ram[14087] = 8'h00;
    ff_ram[14088] = 8'h00;
    ff_ram[14089] = 8'h00;
    ff_ram[14090] = 8'h00;
    ff_ram[14091] = 8'h00;
    ff_ram[14092] = 8'h00;
    ff_ram[14093] = 8'h00;
    ff_ram[14094] = 8'h00;
    ff_ram[14095] = 8'h00;
    ff_ram[14096] = 8'h00;
    ff_ram[14097] = 8'h00;
    ff_ram[14098] = 8'h00;
    ff_ram[14099] = 8'h00;
    ff_ram[14100] = 8'h00;
    ff_ram[14101] = 8'h00;
    ff_ram[14102] = 8'h00;
    ff_ram[14103] = 8'h00;
    ff_ram[14104] = 8'h00;
    ff_ram[14105] = 8'h00;
    ff_ram[14106] = 8'h00;
    ff_ram[14107] = 8'h00;
    ff_ram[14108] = 8'h00;
    ff_ram[14109] = 8'h00;
    ff_ram[14110] = 8'h00;
    ff_ram[14111] = 8'h00;
    ff_ram[14112] = 8'h00;
    ff_ram[14113] = 8'h00;
    ff_ram[14114] = 8'h00;
    ff_ram[14115] = 8'h00;
    ff_ram[14116] = 8'h00;
    ff_ram[14117] = 8'h00;
    ff_ram[14118] = 8'h00;
    ff_ram[14119] = 8'h00;
    ff_ram[14120] = 8'h00;
    ff_ram[14121] = 8'h00;
    ff_ram[14122] = 8'h00;
    ff_ram[14123] = 8'h00;
    ff_ram[14124] = 8'h00;
    ff_ram[14125] = 8'h00;
    ff_ram[14126] = 8'h00;
    ff_ram[14127] = 8'h00;
    ff_ram[14128] = 8'h00;
    ff_ram[14129] = 8'h00;
    ff_ram[14130] = 8'h00;
    ff_ram[14131] = 8'h00;
    ff_ram[14132] = 8'h00;
    ff_ram[14133] = 8'h00;
    ff_ram[14134] = 8'h00;
    ff_ram[14135] = 8'h00;
    ff_ram[14136] = 8'h00;
    ff_ram[14137] = 8'h00;
    ff_ram[14138] = 8'h00;
    ff_ram[14139] = 8'h00;
    ff_ram[14140] = 8'h00;
    ff_ram[14141] = 8'h00;
    ff_ram[14142] = 8'h00;
    ff_ram[14143] = 8'h00;
    ff_ram[14144] = 8'h00;
    ff_ram[14145] = 8'h00;
    ff_ram[14146] = 8'h00;
    ff_ram[14147] = 8'h00;
    ff_ram[14148] = 8'h00;
    ff_ram[14149] = 8'h00;
    ff_ram[14150] = 8'h00;
    ff_ram[14151] = 8'h00;
    ff_ram[14152] = 8'h00;
    ff_ram[14153] = 8'h00;
    ff_ram[14154] = 8'h00;
    ff_ram[14155] = 8'h00;
    ff_ram[14156] = 8'h00;
    ff_ram[14157] = 8'h00;
    ff_ram[14158] = 8'h00;
    ff_ram[14159] = 8'h00;
    ff_ram[14160] = 8'h00;
    ff_ram[14161] = 8'h00;
    ff_ram[14162] = 8'h00;
    ff_ram[14163] = 8'h00;
    ff_ram[14164] = 8'h00;
    ff_ram[14165] = 8'h00;
    ff_ram[14166] = 8'h00;
    ff_ram[14167] = 8'h00;
    ff_ram[14168] = 8'h00;
    ff_ram[14169] = 8'h00;
    ff_ram[14170] = 8'h00;
    ff_ram[14171] = 8'h00;
    ff_ram[14172] = 8'h00;
    ff_ram[14173] = 8'h00;
    ff_ram[14174] = 8'h00;
    ff_ram[14175] = 8'h00;
    ff_ram[14176] = 8'h00;
    ff_ram[14177] = 8'h00;
    ff_ram[14178] = 8'h00;
    ff_ram[14179] = 8'h00;
    ff_ram[14180] = 8'h00;
    ff_ram[14181] = 8'h00;
    ff_ram[14182] = 8'h00;
    ff_ram[14183] = 8'h00;
    ff_ram[14184] = 8'h00;
    ff_ram[14185] = 8'h00;
    ff_ram[14186] = 8'h00;
    ff_ram[14187] = 8'h00;
    ff_ram[14188] = 8'h00;
    ff_ram[14189] = 8'h00;
    ff_ram[14190] = 8'h00;
    ff_ram[14191] = 8'h00;
    ff_ram[14192] = 8'h00;
    ff_ram[14193] = 8'h00;
    ff_ram[14194] = 8'h00;
    ff_ram[14195] = 8'h00;
    ff_ram[14196] = 8'h00;
    ff_ram[14197] = 8'h00;
    ff_ram[14198] = 8'h00;
    ff_ram[14199] = 8'h00;
    ff_ram[14200] = 8'h00;
    ff_ram[14201] = 8'h00;
    ff_ram[14202] = 8'h00;
    ff_ram[14203] = 8'h00;
    ff_ram[14204] = 8'h00;
    ff_ram[14205] = 8'h00;
    ff_ram[14206] = 8'h00;
    ff_ram[14207] = 8'h00;
    ff_ram[14208] = 8'h00;
    ff_ram[14209] = 8'h00;
    ff_ram[14210] = 8'h00;
    ff_ram[14211] = 8'h00;
    ff_ram[14212] = 8'h00;
    ff_ram[14213] = 8'h00;
    ff_ram[14214] = 8'h00;
    ff_ram[14215] = 8'h00;
    ff_ram[14216] = 8'h00;
    ff_ram[14217] = 8'h00;
    ff_ram[14218] = 8'h00;
    ff_ram[14219] = 8'h00;
    ff_ram[14220] = 8'h00;
    ff_ram[14221] = 8'h00;
    ff_ram[14222] = 8'h00;
    ff_ram[14223] = 8'h00;
    ff_ram[14224] = 8'h00;
    ff_ram[14225] = 8'h00;
    ff_ram[14226] = 8'h00;
    ff_ram[14227] = 8'h00;
    ff_ram[14228] = 8'h00;
    ff_ram[14229] = 8'h00;
    ff_ram[14230] = 8'h00;
    ff_ram[14231] = 8'h00;
    ff_ram[14232] = 8'h00;
    ff_ram[14233] = 8'h00;
    ff_ram[14234] = 8'h00;
    ff_ram[14235] = 8'h00;
    ff_ram[14236] = 8'h00;
    ff_ram[14237] = 8'h00;
    ff_ram[14238] = 8'h00;
    ff_ram[14239] = 8'h00;
    ff_ram[14240] = 8'h00;
    ff_ram[14241] = 8'h00;
    ff_ram[14242] = 8'h00;
    ff_ram[14243] = 8'h00;
    ff_ram[14244] = 8'h00;
    ff_ram[14245] = 8'h00;
    ff_ram[14246] = 8'h00;
    ff_ram[14247] = 8'h00;
    ff_ram[14248] = 8'h00;
    ff_ram[14249] = 8'h00;
    ff_ram[14250] = 8'h00;
    ff_ram[14251] = 8'h00;
    ff_ram[14252] = 8'h00;
    ff_ram[14253] = 8'h00;
    ff_ram[14254] = 8'h00;
    ff_ram[14255] = 8'h00;
    ff_ram[14256] = 8'h00;
    ff_ram[14257] = 8'h00;
    ff_ram[14258] = 8'h00;
    ff_ram[14259] = 8'h00;
    ff_ram[14260] = 8'h00;
    ff_ram[14261] = 8'h00;
    ff_ram[14262] = 8'h00;
    ff_ram[14263] = 8'h00;
    ff_ram[14264] = 8'h00;
    ff_ram[14265] = 8'h00;
    ff_ram[14266] = 8'h00;
    ff_ram[14267] = 8'h00;
    ff_ram[14268] = 8'h00;
    ff_ram[14269] = 8'h00;
    ff_ram[14270] = 8'h00;
    ff_ram[14271] = 8'h00;
    ff_ram[14272] = 8'h00;
    ff_ram[14273] = 8'h00;
    ff_ram[14274] = 8'h00;
    ff_ram[14275] = 8'h00;
    ff_ram[14276] = 8'h00;
    ff_ram[14277] = 8'h00;
    ff_ram[14278] = 8'h00;
    ff_ram[14279] = 8'h00;
    ff_ram[14280] = 8'h00;
    ff_ram[14281] = 8'h00;
    ff_ram[14282] = 8'h00;
    ff_ram[14283] = 8'h00;
    ff_ram[14284] = 8'h00;
    ff_ram[14285] = 8'h00;
    ff_ram[14286] = 8'h00;
    ff_ram[14287] = 8'h00;
    ff_ram[14288] = 8'h00;
    ff_ram[14289] = 8'h00;
    ff_ram[14290] = 8'h00;
    ff_ram[14291] = 8'h00;
    ff_ram[14292] = 8'h00;
    ff_ram[14293] = 8'h00;
    ff_ram[14294] = 8'h00;
    ff_ram[14295] = 8'h00;
    ff_ram[14296] = 8'h00;
    ff_ram[14297] = 8'h00;
    ff_ram[14298] = 8'h00;
    ff_ram[14299] = 8'h00;
    ff_ram[14300] = 8'h00;
    ff_ram[14301] = 8'h00;
    ff_ram[14302] = 8'h00;
    ff_ram[14303] = 8'h00;
    ff_ram[14304] = 8'h00;
    ff_ram[14305] = 8'h00;
    ff_ram[14306] = 8'h00;
    ff_ram[14307] = 8'h00;
    ff_ram[14308] = 8'h00;
    ff_ram[14309] = 8'h00;
    ff_ram[14310] = 8'h00;
    ff_ram[14311] = 8'h00;
    ff_ram[14312] = 8'h00;
    ff_ram[14313] = 8'h00;
    ff_ram[14314] = 8'h00;
    ff_ram[14315] = 8'h00;
    ff_ram[14316] = 8'h00;
    ff_ram[14317] = 8'h00;
    ff_ram[14318] = 8'h00;
    ff_ram[14319] = 8'h00;
    ff_ram[14320] = 8'h00;
    ff_ram[14321] = 8'h00;
    ff_ram[14322] = 8'h00;
    ff_ram[14323] = 8'h00;
    ff_ram[14324] = 8'h00;
    ff_ram[14325] = 8'h00;
    ff_ram[14326] = 8'h00;
    ff_ram[14327] = 8'h00;
    ff_ram[14328] = 8'h00;
    ff_ram[14329] = 8'h00;
    ff_ram[14330] = 8'h00;
    ff_ram[14331] = 8'h00;
    ff_ram[14332] = 8'h00;
    ff_ram[14333] = 8'h00;
    ff_ram[14334] = 8'h00;
    ff_ram[14335] = 8'h00;
    ff_ram[14336] = 8'h00;
    ff_ram[14337] = 8'h00;
    ff_ram[14338] = 8'h00;
    ff_ram[14339] = 8'h00;
    ff_ram[14340] = 8'h00;
    ff_ram[14341] = 8'h00;
    ff_ram[14342] = 8'h00;
    ff_ram[14343] = 8'h00;
    ff_ram[14344] = 8'h00;
    ff_ram[14345] = 8'h00;
    ff_ram[14346] = 8'h00;
    ff_ram[14347] = 8'h00;
    ff_ram[14348] = 8'h00;
    ff_ram[14349] = 8'h00;
    ff_ram[14350] = 8'h00;
    ff_ram[14351] = 8'h00;
    ff_ram[14352] = 8'h00;
    ff_ram[14353] = 8'h00;
    ff_ram[14354] = 8'h00;
    ff_ram[14355] = 8'h00;
    ff_ram[14356] = 8'h00;
    ff_ram[14357] = 8'h00;
    ff_ram[14358] = 8'h00;
    ff_ram[14359] = 8'h00;
    ff_ram[14360] = 8'h00;
    ff_ram[14361] = 8'h00;
    ff_ram[14362] = 8'h00;
    ff_ram[14363] = 8'h00;
    ff_ram[14364] = 8'h00;
    ff_ram[14365] = 8'h00;
    ff_ram[14366] = 8'h00;
    ff_ram[14367] = 8'h00;
    ff_ram[14368] = 8'h00;
    ff_ram[14369] = 8'h00;
    ff_ram[14370] = 8'h00;
    ff_ram[14371] = 8'h00;
    ff_ram[14372] = 8'h00;
    ff_ram[14373] = 8'h00;
    ff_ram[14374] = 8'h00;
    ff_ram[14375] = 8'h00;
    ff_ram[14376] = 8'h00;
    ff_ram[14377] = 8'h00;
    ff_ram[14378] = 8'h00;
    ff_ram[14379] = 8'h00;
    ff_ram[14380] = 8'h00;
    ff_ram[14381] = 8'h00;
    ff_ram[14382] = 8'h00;
    ff_ram[14383] = 8'h00;
    ff_ram[14384] = 8'h00;
    ff_ram[14385] = 8'h00;
    ff_ram[14386] = 8'h00;
    ff_ram[14387] = 8'h00;
    ff_ram[14388] = 8'h00;
    ff_ram[14389] = 8'h00;
    ff_ram[14390] = 8'h00;
    ff_ram[14391] = 8'h00;
    ff_ram[14392] = 8'h00;
    ff_ram[14393] = 8'h00;
    ff_ram[14394] = 8'h00;
    ff_ram[14395] = 8'h00;
    ff_ram[14396] = 8'h00;
    ff_ram[14397] = 8'h00;
    ff_ram[14398] = 8'h00;
    ff_ram[14399] = 8'h00;
    ff_ram[14400] = 8'h00;
    ff_ram[14401] = 8'h00;
    ff_ram[14402] = 8'h00;
    ff_ram[14403] = 8'h00;
    ff_ram[14404] = 8'h00;
    ff_ram[14405] = 8'h00;
    ff_ram[14406] = 8'h00;
    ff_ram[14407] = 8'h00;
    ff_ram[14408] = 8'h00;
    ff_ram[14409] = 8'h00;
    ff_ram[14410] = 8'h00;
    ff_ram[14411] = 8'h00;
    ff_ram[14412] = 8'h00;
    ff_ram[14413] = 8'h00;
    ff_ram[14414] = 8'h00;
    ff_ram[14415] = 8'h00;
    ff_ram[14416] = 8'h00;
    ff_ram[14417] = 8'h00;
    ff_ram[14418] = 8'h00;
    ff_ram[14419] = 8'h00;
    ff_ram[14420] = 8'h00;
    ff_ram[14421] = 8'h00;
    ff_ram[14422] = 8'h00;
    ff_ram[14423] = 8'h00;
    ff_ram[14424] = 8'h00;
    ff_ram[14425] = 8'h00;
    ff_ram[14426] = 8'h00;
    ff_ram[14427] = 8'h00;
    ff_ram[14428] = 8'h00;
    ff_ram[14429] = 8'h00;
    ff_ram[14430] = 8'h00;
    ff_ram[14431] = 8'h00;
    ff_ram[14432] = 8'h00;
    ff_ram[14433] = 8'h00;
    ff_ram[14434] = 8'h00;
    ff_ram[14435] = 8'h00;
    ff_ram[14436] = 8'h00;
    ff_ram[14437] = 8'h00;
    ff_ram[14438] = 8'h00;
    ff_ram[14439] = 8'h00;
    ff_ram[14440] = 8'h00;
    ff_ram[14441] = 8'h00;
    ff_ram[14442] = 8'h00;
    ff_ram[14443] = 8'h00;
    ff_ram[14444] = 8'h00;
    ff_ram[14445] = 8'h00;
    ff_ram[14446] = 8'h00;
    ff_ram[14447] = 8'h00;
    ff_ram[14448] = 8'h00;
    ff_ram[14449] = 8'h00;
    ff_ram[14450] = 8'h00;
    ff_ram[14451] = 8'h00;
    ff_ram[14452] = 8'h00;
    ff_ram[14453] = 8'h00;
    ff_ram[14454] = 8'h00;
    ff_ram[14455] = 8'h00;
    ff_ram[14456] = 8'h00;
    ff_ram[14457] = 8'h00;
    ff_ram[14458] = 8'h00;
    ff_ram[14459] = 8'h00;
    ff_ram[14460] = 8'h00;
    ff_ram[14461] = 8'h00;
    ff_ram[14462] = 8'h00;
    ff_ram[14463] = 8'h00;
    ff_ram[14464] = 8'h00;
    ff_ram[14465] = 8'h00;
    ff_ram[14466] = 8'h00;
    ff_ram[14467] = 8'h00;
    ff_ram[14468] = 8'h00;
    ff_ram[14469] = 8'h00;
    ff_ram[14470] = 8'h00;
    ff_ram[14471] = 8'h00;
    ff_ram[14472] = 8'h00;
    ff_ram[14473] = 8'h00;
    ff_ram[14474] = 8'h00;
    ff_ram[14475] = 8'h00;
    ff_ram[14476] = 8'h00;
    ff_ram[14477] = 8'h00;
    ff_ram[14478] = 8'h00;
    ff_ram[14479] = 8'h00;
    ff_ram[14480] = 8'h00;
    ff_ram[14481] = 8'h00;
    ff_ram[14482] = 8'h00;
    ff_ram[14483] = 8'h00;
    ff_ram[14484] = 8'h00;
    ff_ram[14485] = 8'h00;
    ff_ram[14486] = 8'h00;
    ff_ram[14487] = 8'h00;
    ff_ram[14488] = 8'h00;
    ff_ram[14489] = 8'h00;
    ff_ram[14490] = 8'h00;
    ff_ram[14491] = 8'h00;
    ff_ram[14492] = 8'h00;
    ff_ram[14493] = 8'h00;
    ff_ram[14494] = 8'h00;
    ff_ram[14495] = 8'h00;
    ff_ram[14496] = 8'h00;
    ff_ram[14497] = 8'h00;
    ff_ram[14498] = 8'h00;
    ff_ram[14499] = 8'h00;
    ff_ram[14500] = 8'h00;
    ff_ram[14501] = 8'h00;
    ff_ram[14502] = 8'h00;
    ff_ram[14503] = 8'h00;
    ff_ram[14504] = 8'h00;
    ff_ram[14505] = 8'h00;
    ff_ram[14506] = 8'h00;
    ff_ram[14507] = 8'h00;
    ff_ram[14508] = 8'h00;
    ff_ram[14509] = 8'h00;
    ff_ram[14510] = 8'h00;
    ff_ram[14511] = 8'h00;
    ff_ram[14512] = 8'h00;
    ff_ram[14513] = 8'h00;
    ff_ram[14514] = 8'h00;
    ff_ram[14515] = 8'h00;
    ff_ram[14516] = 8'h00;
    ff_ram[14517] = 8'h00;
    ff_ram[14518] = 8'h00;
    ff_ram[14519] = 8'h00;
    ff_ram[14520] = 8'h00;
    ff_ram[14521] = 8'h00;
    ff_ram[14522] = 8'h00;
    ff_ram[14523] = 8'h00;
    ff_ram[14524] = 8'h00;
    ff_ram[14525] = 8'h00;
    ff_ram[14526] = 8'h00;
    ff_ram[14527] = 8'h00;
    ff_ram[14528] = 8'h00;
    ff_ram[14529] = 8'h00;
    ff_ram[14530] = 8'h00;
    ff_ram[14531] = 8'h00;
    ff_ram[14532] = 8'h00;
    ff_ram[14533] = 8'h00;
    ff_ram[14534] = 8'h00;
    ff_ram[14535] = 8'h00;
    ff_ram[14536] = 8'h00;
    ff_ram[14537] = 8'h00;
    ff_ram[14538] = 8'h00;
    ff_ram[14539] = 8'h00;
    ff_ram[14540] = 8'h00;
    ff_ram[14541] = 8'h00;
    ff_ram[14542] = 8'h00;
    ff_ram[14543] = 8'h00;
    ff_ram[14544] = 8'h00;
    ff_ram[14545] = 8'h00;
    ff_ram[14546] = 8'h00;
    ff_ram[14547] = 8'h00;
    ff_ram[14548] = 8'h00;
    ff_ram[14549] = 8'h00;
    ff_ram[14550] = 8'h00;
    ff_ram[14551] = 8'h00;
    ff_ram[14552] = 8'h00;
    ff_ram[14553] = 8'h00;
    ff_ram[14554] = 8'h00;
    ff_ram[14555] = 8'h00;
    ff_ram[14556] = 8'h00;
    ff_ram[14557] = 8'h00;
    ff_ram[14558] = 8'h00;
    ff_ram[14559] = 8'h00;
    ff_ram[14560] = 8'h00;
    ff_ram[14561] = 8'h00;
    ff_ram[14562] = 8'h00;
    ff_ram[14563] = 8'h00;
    ff_ram[14564] = 8'h00;
    ff_ram[14565] = 8'h00;
    ff_ram[14566] = 8'h00;
    ff_ram[14567] = 8'h00;
    ff_ram[14568] = 8'h00;
    ff_ram[14569] = 8'h00;
    ff_ram[14570] = 8'h00;
    ff_ram[14571] = 8'h00;
    ff_ram[14572] = 8'h00;
    ff_ram[14573] = 8'h00;
    ff_ram[14574] = 8'h00;
    ff_ram[14575] = 8'h00;
    ff_ram[14576] = 8'h00;
    ff_ram[14577] = 8'h00;
    ff_ram[14578] = 8'h00;
    ff_ram[14579] = 8'h00;
    ff_ram[14580] = 8'h00;
    ff_ram[14581] = 8'h00;
    ff_ram[14582] = 8'h00;
    ff_ram[14583] = 8'h00;
    ff_ram[14584] = 8'h00;
    ff_ram[14585] = 8'h00;
    ff_ram[14586] = 8'h00;
    ff_ram[14587] = 8'h00;
    ff_ram[14588] = 8'h00;
    ff_ram[14589] = 8'h00;
    ff_ram[14590] = 8'h00;
    ff_ram[14591] = 8'h00;
    ff_ram[14592] = 8'h00;
    ff_ram[14593] = 8'h00;
    ff_ram[14594] = 8'h00;
    ff_ram[14595] = 8'h00;
    ff_ram[14596] = 8'h00;
    ff_ram[14597] = 8'h00;
    ff_ram[14598] = 8'h00;
    ff_ram[14599] = 8'h00;
    ff_ram[14600] = 8'h00;
    ff_ram[14601] = 8'h00;
    ff_ram[14602] = 8'h00;
    ff_ram[14603] = 8'h00;
    ff_ram[14604] = 8'h00;
    ff_ram[14605] = 8'h00;
    ff_ram[14606] = 8'h00;
    ff_ram[14607] = 8'h00;
    ff_ram[14608] = 8'h00;
    ff_ram[14609] = 8'h00;
    ff_ram[14610] = 8'h00;
    ff_ram[14611] = 8'h00;
    ff_ram[14612] = 8'h00;
    ff_ram[14613] = 8'h00;
    ff_ram[14614] = 8'h00;
    ff_ram[14615] = 8'h00;
    ff_ram[14616] = 8'h00;
    ff_ram[14617] = 8'h00;
    ff_ram[14618] = 8'h00;
    ff_ram[14619] = 8'h00;
    ff_ram[14620] = 8'h00;
    ff_ram[14621] = 8'h00;
    ff_ram[14622] = 8'h00;
    ff_ram[14623] = 8'h00;
    ff_ram[14624] = 8'h00;
    ff_ram[14625] = 8'h00;
    ff_ram[14626] = 8'h00;
    ff_ram[14627] = 8'h00;
    ff_ram[14628] = 8'h00;
    ff_ram[14629] = 8'h00;
    ff_ram[14630] = 8'h00;
    ff_ram[14631] = 8'h00;
    ff_ram[14632] = 8'h00;
    ff_ram[14633] = 8'h00;
    ff_ram[14634] = 8'h00;
    ff_ram[14635] = 8'h00;
    ff_ram[14636] = 8'h00;
    ff_ram[14637] = 8'h00;
    ff_ram[14638] = 8'h00;
    ff_ram[14639] = 8'h00;
    ff_ram[14640] = 8'h00;
    ff_ram[14641] = 8'h00;
    ff_ram[14642] = 8'h00;
    ff_ram[14643] = 8'h00;
    ff_ram[14644] = 8'h00;
    ff_ram[14645] = 8'h00;
    ff_ram[14646] = 8'h00;
    ff_ram[14647] = 8'h00;
    ff_ram[14648] = 8'h00;
    ff_ram[14649] = 8'h00;
    ff_ram[14650] = 8'h00;
    ff_ram[14651] = 8'h00;
    ff_ram[14652] = 8'h00;
    ff_ram[14653] = 8'h00;
    ff_ram[14654] = 8'h00;
    ff_ram[14655] = 8'h00;
    ff_ram[14656] = 8'h00;
    ff_ram[14657] = 8'h00;
    ff_ram[14658] = 8'h00;
    ff_ram[14659] = 8'h00;
    ff_ram[14660] = 8'h00;
    ff_ram[14661] = 8'h00;
    ff_ram[14662] = 8'h00;
    ff_ram[14663] = 8'h00;
    ff_ram[14664] = 8'h00;
    ff_ram[14665] = 8'h00;
    ff_ram[14666] = 8'h00;
    ff_ram[14667] = 8'h00;
    ff_ram[14668] = 8'h00;
    ff_ram[14669] = 8'h00;
    ff_ram[14670] = 8'h00;
    ff_ram[14671] = 8'h00;
    ff_ram[14672] = 8'h00;
    ff_ram[14673] = 8'h00;
    ff_ram[14674] = 8'h00;
    ff_ram[14675] = 8'h00;
    ff_ram[14676] = 8'h00;
    ff_ram[14677] = 8'h00;
    ff_ram[14678] = 8'h00;
    ff_ram[14679] = 8'h00;
    ff_ram[14680] = 8'h00;
    ff_ram[14681] = 8'h00;
    ff_ram[14682] = 8'h00;
    ff_ram[14683] = 8'h00;
    ff_ram[14684] = 8'h00;
    ff_ram[14685] = 8'h00;
    ff_ram[14686] = 8'h00;
    ff_ram[14687] = 8'h00;
    ff_ram[14688] = 8'h00;
    ff_ram[14689] = 8'h00;
    ff_ram[14690] = 8'h00;
    ff_ram[14691] = 8'h00;
    ff_ram[14692] = 8'h00;
    ff_ram[14693] = 8'h00;
    ff_ram[14694] = 8'h00;
    ff_ram[14695] = 8'h00;
    ff_ram[14696] = 8'h00;
    ff_ram[14697] = 8'h00;
    ff_ram[14698] = 8'h00;
    ff_ram[14699] = 8'h00;
    ff_ram[14700] = 8'h00;
    ff_ram[14701] = 8'h00;
    ff_ram[14702] = 8'h00;
    ff_ram[14703] = 8'h00;
    ff_ram[14704] = 8'h00;
    ff_ram[14705] = 8'h00;
    ff_ram[14706] = 8'h00;
    ff_ram[14707] = 8'h00;
    ff_ram[14708] = 8'h00;
    ff_ram[14709] = 8'h00;
    ff_ram[14710] = 8'h00;
    ff_ram[14711] = 8'h00;
    ff_ram[14712] = 8'h00;
    ff_ram[14713] = 8'h00;
    ff_ram[14714] = 8'h00;
    ff_ram[14715] = 8'h00;
    ff_ram[14716] = 8'h00;
    ff_ram[14717] = 8'h00;
    ff_ram[14718] = 8'h00;
    ff_ram[14719] = 8'h00;
    ff_ram[14720] = 8'h00;
    ff_ram[14721] = 8'h00;
    ff_ram[14722] = 8'h00;
    ff_ram[14723] = 8'h00;
    ff_ram[14724] = 8'h00;
    ff_ram[14725] = 8'h00;
    ff_ram[14726] = 8'h00;
    ff_ram[14727] = 8'h00;
    ff_ram[14728] = 8'h00;
    ff_ram[14729] = 8'h00;
    ff_ram[14730] = 8'h00;
    ff_ram[14731] = 8'h00;
    ff_ram[14732] = 8'h00;
    ff_ram[14733] = 8'h00;
    ff_ram[14734] = 8'h00;
    ff_ram[14735] = 8'h00;
    ff_ram[14736] = 8'h00;
    ff_ram[14737] = 8'h00;
    ff_ram[14738] = 8'h00;
    ff_ram[14739] = 8'h00;
    ff_ram[14740] = 8'h00;
    ff_ram[14741] = 8'h00;
    ff_ram[14742] = 8'h00;
    ff_ram[14743] = 8'h00;
    ff_ram[14744] = 8'h00;
    ff_ram[14745] = 8'h00;
    ff_ram[14746] = 8'h00;
    ff_ram[14747] = 8'h00;
    ff_ram[14748] = 8'h00;
    ff_ram[14749] = 8'h00;
    ff_ram[14750] = 8'h00;
    ff_ram[14751] = 8'h00;
    ff_ram[14752] = 8'h00;
    ff_ram[14753] = 8'h00;
    ff_ram[14754] = 8'h00;
    ff_ram[14755] = 8'h00;
    ff_ram[14756] = 8'h00;
    ff_ram[14757] = 8'h00;
    ff_ram[14758] = 8'h00;
    ff_ram[14759] = 8'h00;
    ff_ram[14760] = 8'h00;
    ff_ram[14761] = 8'h00;
    ff_ram[14762] = 8'h00;
    ff_ram[14763] = 8'h00;
    ff_ram[14764] = 8'h00;
    ff_ram[14765] = 8'h00;
    ff_ram[14766] = 8'h00;
    ff_ram[14767] = 8'h00;
    ff_ram[14768] = 8'h00;
    ff_ram[14769] = 8'h00;
    ff_ram[14770] = 8'h00;
    ff_ram[14771] = 8'h00;
    ff_ram[14772] = 8'h00;
    ff_ram[14773] = 8'h00;
    ff_ram[14774] = 8'h00;
    ff_ram[14775] = 8'h00;
    ff_ram[14776] = 8'h00;
    ff_ram[14777] = 8'h00;
    ff_ram[14778] = 8'h00;
    ff_ram[14779] = 8'h00;
    ff_ram[14780] = 8'h00;
    ff_ram[14781] = 8'h00;
    ff_ram[14782] = 8'h00;
    ff_ram[14783] = 8'h00;
    ff_ram[14784] = 8'h00;
    ff_ram[14785] = 8'h00;
    ff_ram[14786] = 8'h00;
    ff_ram[14787] = 8'h00;
    ff_ram[14788] = 8'h00;
    ff_ram[14789] = 8'h00;
    ff_ram[14790] = 8'h00;
    ff_ram[14791] = 8'h00;
    ff_ram[14792] = 8'h00;
    ff_ram[14793] = 8'h00;
    ff_ram[14794] = 8'h00;
    ff_ram[14795] = 8'h00;
    ff_ram[14796] = 8'h00;
    ff_ram[14797] = 8'h00;
    ff_ram[14798] = 8'h00;
    ff_ram[14799] = 8'h00;
    ff_ram[14800] = 8'h00;
    ff_ram[14801] = 8'h00;
    ff_ram[14802] = 8'h00;
    ff_ram[14803] = 8'h00;
    ff_ram[14804] = 8'h00;
    ff_ram[14805] = 8'h00;
    ff_ram[14806] = 8'h00;
    ff_ram[14807] = 8'h00;
    ff_ram[14808] = 8'h00;
    ff_ram[14809] = 8'h00;
    ff_ram[14810] = 8'h00;
    ff_ram[14811] = 8'h00;
    ff_ram[14812] = 8'h00;
    ff_ram[14813] = 8'h00;
    ff_ram[14814] = 8'h00;
    ff_ram[14815] = 8'h00;
    ff_ram[14816] = 8'h00;
    ff_ram[14817] = 8'h00;
    ff_ram[14818] = 8'h00;
    ff_ram[14819] = 8'h00;
    ff_ram[14820] = 8'h00;
    ff_ram[14821] = 8'h00;
    ff_ram[14822] = 8'h00;
    ff_ram[14823] = 8'h00;
    ff_ram[14824] = 8'h00;
    ff_ram[14825] = 8'h00;
    ff_ram[14826] = 8'h00;
    ff_ram[14827] = 8'h00;
    ff_ram[14828] = 8'h00;
    ff_ram[14829] = 8'h00;
    ff_ram[14830] = 8'h00;
    ff_ram[14831] = 8'h00;
    ff_ram[14832] = 8'h00;
    ff_ram[14833] = 8'h00;
    ff_ram[14834] = 8'h00;
    ff_ram[14835] = 8'h00;
    ff_ram[14836] = 8'h00;
    ff_ram[14837] = 8'h00;
    ff_ram[14838] = 8'h00;
    ff_ram[14839] = 8'h00;
    ff_ram[14840] = 8'h00;
    ff_ram[14841] = 8'h00;
    ff_ram[14842] = 8'h00;
    ff_ram[14843] = 8'h00;
    ff_ram[14844] = 8'h00;
    ff_ram[14845] = 8'h00;
    ff_ram[14846] = 8'h00;
    ff_ram[14847] = 8'h00;
    ff_ram[14848] = 8'h00;
    ff_ram[14849] = 8'h00;
    ff_ram[14850] = 8'h00;
    ff_ram[14851] = 8'h00;
    ff_ram[14852] = 8'h00;
    ff_ram[14853] = 8'h00;
    ff_ram[14854] = 8'h00;
    ff_ram[14855] = 8'h00;
    ff_ram[14856] = 8'h00;
    ff_ram[14857] = 8'h00;
    ff_ram[14858] = 8'h00;
    ff_ram[14859] = 8'h00;
    ff_ram[14860] = 8'h00;
    ff_ram[14861] = 8'h00;
    ff_ram[14862] = 8'h00;
    ff_ram[14863] = 8'h00;
    ff_ram[14864] = 8'h00;
    ff_ram[14865] = 8'h00;
    ff_ram[14866] = 8'h00;
    ff_ram[14867] = 8'h00;
    ff_ram[14868] = 8'h00;
    ff_ram[14869] = 8'h00;
    ff_ram[14870] = 8'h00;
    ff_ram[14871] = 8'h00;
    ff_ram[14872] = 8'h00;
    ff_ram[14873] = 8'h00;
    ff_ram[14874] = 8'h00;
    ff_ram[14875] = 8'h00;
    ff_ram[14876] = 8'h00;
    ff_ram[14877] = 8'h00;
    ff_ram[14878] = 8'h00;
    ff_ram[14879] = 8'h00;
    ff_ram[14880] = 8'h00;
    ff_ram[14881] = 8'h00;
    ff_ram[14882] = 8'h00;
    ff_ram[14883] = 8'h00;
    ff_ram[14884] = 8'h00;
    ff_ram[14885] = 8'h00;
    ff_ram[14886] = 8'h00;
    ff_ram[14887] = 8'h00;
    ff_ram[14888] = 8'h00;
    ff_ram[14889] = 8'h00;
    ff_ram[14890] = 8'h00;
    ff_ram[14891] = 8'h00;
    ff_ram[14892] = 8'h00;
    ff_ram[14893] = 8'h00;
    ff_ram[14894] = 8'h00;
    ff_ram[14895] = 8'h00;
    ff_ram[14896] = 8'h00;
    ff_ram[14897] = 8'h00;
    ff_ram[14898] = 8'h00;
    ff_ram[14899] = 8'h00;
    ff_ram[14900] = 8'h00;
    ff_ram[14901] = 8'h00;
    ff_ram[14902] = 8'h00;
    ff_ram[14903] = 8'h00;
    ff_ram[14904] = 8'h00;
    ff_ram[14905] = 8'h00;
    ff_ram[14906] = 8'h00;
    ff_ram[14907] = 8'h00;
    ff_ram[14908] = 8'h00;
    ff_ram[14909] = 8'h00;
    ff_ram[14910] = 8'h00;
    ff_ram[14911] = 8'h00;
    ff_ram[14912] = 8'h00;
    ff_ram[14913] = 8'h00;
    ff_ram[14914] = 8'h00;
    ff_ram[14915] = 8'h00;
    ff_ram[14916] = 8'h00;
    ff_ram[14917] = 8'h00;
    ff_ram[14918] = 8'h00;
    ff_ram[14919] = 8'h00;
    ff_ram[14920] = 8'h00;
    ff_ram[14921] = 8'h00;
    ff_ram[14922] = 8'h00;
    ff_ram[14923] = 8'h00;
    ff_ram[14924] = 8'h00;
    ff_ram[14925] = 8'h00;
    ff_ram[14926] = 8'h00;
    ff_ram[14927] = 8'h00;
    ff_ram[14928] = 8'h00;
    ff_ram[14929] = 8'h00;
    ff_ram[14930] = 8'h00;
    ff_ram[14931] = 8'h00;
    ff_ram[14932] = 8'h00;
    ff_ram[14933] = 8'h00;
    ff_ram[14934] = 8'h00;
    ff_ram[14935] = 8'h00;
    ff_ram[14936] = 8'h00;
    ff_ram[14937] = 8'h00;
    ff_ram[14938] = 8'h00;
    ff_ram[14939] = 8'h00;
    ff_ram[14940] = 8'h00;
    ff_ram[14941] = 8'h00;
    ff_ram[14942] = 8'h00;
    ff_ram[14943] = 8'h00;
    ff_ram[14944] = 8'h00;
    ff_ram[14945] = 8'h00;
    ff_ram[14946] = 8'h00;
    ff_ram[14947] = 8'h00;
    ff_ram[14948] = 8'h00;
    ff_ram[14949] = 8'h00;
    ff_ram[14950] = 8'h00;
    ff_ram[14951] = 8'h00;
    ff_ram[14952] = 8'h00;
    ff_ram[14953] = 8'h00;
    ff_ram[14954] = 8'h00;
    ff_ram[14955] = 8'h00;
    ff_ram[14956] = 8'h00;
    ff_ram[14957] = 8'h00;
    ff_ram[14958] = 8'h00;
    ff_ram[14959] = 8'h00;
    ff_ram[14960] = 8'h00;
    ff_ram[14961] = 8'h00;
    ff_ram[14962] = 8'h00;
    ff_ram[14963] = 8'h00;
    ff_ram[14964] = 8'h00;
    ff_ram[14965] = 8'h00;
    ff_ram[14966] = 8'h00;
    ff_ram[14967] = 8'h00;
    ff_ram[14968] = 8'h00;
    ff_ram[14969] = 8'h00;
    ff_ram[14970] = 8'h00;
    ff_ram[14971] = 8'h00;
    ff_ram[14972] = 8'h00;
    ff_ram[14973] = 8'h00;
    ff_ram[14974] = 8'h00;
    ff_ram[14975] = 8'h00;
    ff_ram[14976] = 8'h00;
    ff_ram[14977] = 8'h00;
    ff_ram[14978] = 8'h00;
    ff_ram[14979] = 8'h00;
    ff_ram[14980] = 8'h00;
    ff_ram[14981] = 8'h00;
    ff_ram[14982] = 8'h00;
    ff_ram[14983] = 8'h00;
    ff_ram[14984] = 8'h00;
    ff_ram[14985] = 8'h00;
    ff_ram[14986] = 8'h00;
    ff_ram[14987] = 8'h00;
    ff_ram[14988] = 8'h00;
    ff_ram[14989] = 8'h00;
    ff_ram[14990] = 8'h00;
    ff_ram[14991] = 8'h00;
    ff_ram[14992] = 8'h00;
    ff_ram[14993] = 8'h00;
    ff_ram[14994] = 8'h00;
    ff_ram[14995] = 8'h00;
    ff_ram[14996] = 8'h00;
    ff_ram[14997] = 8'h00;
    ff_ram[14998] = 8'h00;
    ff_ram[14999] = 8'h00;
    ff_ram[15000] = 8'h00;
    ff_ram[15001] = 8'h00;
    ff_ram[15002] = 8'h00;
    ff_ram[15003] = 8'h00;
    ff_ram[15004] = 8'h00;
    ff_ram[15005] = 8'h00;
    ff_ram[15006] = 8'h00;
    ff_ram[15007] = 8'h00;
    ff_ram[15008] = 8'h00;
    ff_ram[15009] = 8'h00;
    ff_ram[15010] = 8'h00;
    ff_ram[15011] = 8'h00;
    ff_ram[15012] = 8'h00;
    ff_ram[15013] = 8'h00;
    ff_ram[15014] = 8'h00;
    ff_ram[15015] = 8'h00;
    ff_ram[15016] = 8'h00;
    ff_ram[15017] = 8'h00;
    ff_ram[15018] = 8'h00;
    ff_ram[15019] = 8'h00;
    ff_ram[15020] = 8'h00;
    ff_ram[15021] = 8'h00;
    ff_ram[15022] = 8'h00;
    ff_ram[15023] = 8'h00;
    ff_ram[15024] = 8'h00;
    ff_ram[15025] = 8'h00;
    ff_ram[15026] = 8'h00;
    ff_ram[15027] = 8'h00;
    ff_ram[15028] = 8'h00;
    ff_ram[15029] = 8'h00;
    ff_ram[15030] = 8'h00;
    ff_ram[15031] = 8'h00;
    ff_ram[15032] = 8'h00;
    ff_ram[15033] = 8'h00;
    ff_ram[15034] = 8'h00;
    ff_ram[15035] = 8'h00;
    ff_ram[15036] = 8'h00;
    ff_ram[15037] = 8'h00;
    ff_ram[15038] = 8'h00;
    ff_ram[15039] = 8'h00;
    ff_ram[15040] = 8'h00;
    ff_ram[15041] = 8'h00;
    ff_ram[15042] = 8'h00;
    ff_ram[15043] = 8'h00;
    ff_ram[15044] = 8'h00;
    ff_ram[15045] = 8'h00;
    ff_ram[15046] = 8'h00;
    ff_ram[15047] = 8'h00;
    ff_ram[15048] = 8'h00;
    ff_ram[15049] = 8'h00;
    ff_ram[15050] = 8'h00;
    ff_ram[15051] = 8'h00;
    ff_ram[15052] = 8'h00;
    ff_ram[15053] = 8'h00;
    ff_ram[15054] = 8'h00;
    ff_ram[15055] = 8'h00;
    ff_ram[15056] = 8'h00;
    ff_ram[15057] = 8'h00;
    ff_ram[15058] = 8'h00;
    ff_ram[15059] = 8'h00;
    ff_ram[15060] = 8'h00;
    ff_ram[15061] = 8'h00;
    ff_ram[15062] = 8'h00;
    ff_ram[15063] = 8'h00;
    ff_ram[15064] = 8'h00;
    ff_ram[15065] = 8'h00;
    ff_ram[15066] = 8'h00;
    ff_ram[15067] = 8'h00;
    ff_ram[15068] = 8'h00;
    ff_ram[15069] = 8'h00;
    ff_ram[15070] = 8'h00;
    ff_ram[15071] = 8'h00;
    ff_ram[15072] = 8'h00;
    ff_ram[15073] = 8'h00;
    ff_ram[15074] = 8'h00;
    ff_ram[15075] = 8'h00;
    ff_ram[15076] = 8'h00;
    ff_ram[15077] = 8'h00;
    ff_ram[15078] = 8'h00;
    ff_ram[15079] = 8'h00;
    ff_ram[15080] = 8'h00;
    ff_ram[15081] = 8'h00;
    ff_ram[15082] = 8'h00;
    ff_ram[15083] = 8'h00;
    ff_ram[15084] = 8'h00;
    ff_ram[15085] = 8'h00;
    ff_ram[15086] = 8'h00;
    ff_ram[15087] = 8'h00;
    ff_ram[15088] = 8'h00;
    ff_ram[15089] = 8'h00;
    ff_ram[15090] = 8'h00;
    ff_ram[15091] = 8'h00;
    ff_ram[15092] = 8'h00;
    ff_ram[15093] = 8'h00;
    ff_ram[15094] = 8'h00;
    ff_ram[15095] = 8'h00;
    ff_ram[15096] = 8'h00;
    ff_ram[15097] = 8'h00;
    ff_ram[15098] = 8'h00;
    ff_ram[15099] = 8'h00;
    ff_ram[15100] = 8'h00;
    ff_ram[15101] = 8'h00;
    ff_ram[15102] = 8'h00;
    ff_ram[15103] = 8'h00;
    ff_ram[15104] = 8'h00;
    ff_ram[15105] = 8'h00;
    ff_ram[15106] = 8'h00;
    ff_ram[15107] = 8'h00;
    ff_ram[15108] = 8'h00;
    ff_ram[15109] = 8'h00;
    ff_ram[15110] = 8'h00;
    ff_ram[15111] = 8'h00;
    ff_ram[15112] = 8'h00;
    ff_ram[15113] = 8'h00;
    ff_ram[15114] = 8'h00;
    ff_ram[15115] = 8'h00;
    ff_ram[15116] = 8'h00;
    ff_ram[15117] = 8'h00;
    ff_ram[15118] = 8'h00;
    ff_ram[15119] = 8'h00;
    ff_ram[15120] = 8'h00;
    ff_ram[15121] = 8'h00;
    ff_ram[15122] = 8'h00;
    ff_ram[15123] = 8'h00;
    ff_ram[15124] = 8'h00;
    ff_ram[15125] = 8'h00;
    ff_ram[15126] = 8'h00;
    ff_ram[15127] = 8'h00;
    ff_ram[15128] = 8'h00;
    ff_ram[15129] = 8'h00;
    ff_ram[15130] = 8'h00;
    ff_ram[15131] = 8'h00;
    ff_ram[15132] = 8'h00;
    ff_ram[15133] = 8'h00;
    ff_ram[15134] = 8'h00;
    ff_ram[15135] = 8'h00;
    ff_ram[15136] = 8'h00;
    ff_ram[15137] = 8'h00;
    ff_ram[15138] = 8'h00;
    ff_ram[15139] = 8'h00;
    ff_ram[15140] = 8'h00;
    ff_ram[15141] = 8'h00;
    ff_ram[15142] = 8'h00;
    ff_ram[15143] = 8'h00;
    ff_ram[15144] = 8'h00;
    ff_ram[15145] = 8'h00;
    ff_ram[15146] = 8'h00;
    ff_ram[15147] = 8'h00;
    ff_ram[15148] = 8'h00;
    ff_ram[15149] = 8'h00;
    ff_ram[15150] = 8'h00;
    ff_ram[15151] = 8'h00;
    ff_ram[15152] = 8'h00;
    ff_ram[15153] = 8'h00;
    ff_ram[15154] = 8'h00;
    ff_ram[15155] = 8'h00;
    ff_ram[15156] = 8'h00;
    ff_ram[15157] = 8'h00;
    ff_ram[15158] = 8'h00;
    ff_ram[15159] = 8'h00;
    ff_ram[15160] = 8'h00;
    ff_ram[15161] = 8'h00;
    ff_ram[15162] = 8'h00;
    ff_ram[15163] = 8'h00;
    ff_ram[15164] = 8'h00;
    ff_ram[15165] = 8'h00;
    ff_ram[15166] = 8'h00;
    ff_ram[15167] = 8'h00;
    ff_ram[15168] = 8'h00;
    ff_ram[15169] = 8'h00;
    ff_ram[15170] = 8'h00;
    ff_ram[15171] = 8'h00;
    ff_ram[15172] = 8'h00;
    ff_ram[15173] = 8'h00;
    ff_ram[15174] = 8'h00;
    ff_ram[15175] = 8'h00;
    ff_ram[15176] = 8'h00;
    ff_ram[15177] = 8'h00;
    ff_ram[15178] = 8'h00;
    ff_ram[15179] = 8'h00;
    ff_ram[15180] = 8'h00;
    ff_ram[15181] = 8'h00;
    ff_ram[15182] = 8'h00;
    ff_ram[15183] = 8'h00;
    ff_ram[15184] = 8'h00;
    ff_ram[15185] = 8'h00;
    ff_ram[15186] = 8'h00;
    ff_ram[15187] = 8'h00;
    ff_ram[15188] = 8'h00;
    ff_ram[15189] = 8'h00;
    ff_ram[15190] = 8'h00;
    ff_ram[15191] = 8'h00;
    ff_ram[15192] = 8'h00;
    ff_ram[15193] = 8'h00;
    ff_ram[15194] = 8'h00;
    ff_ram[15195] = 8'h00;
    ff_ram[15196] = 8'h00;
    ff_ram[15197] = 8'h00;
    ff_ram[15198] = 8'h00;
    ff_ram[15199] = 8'h00;
    ff_ram[15200] = 8'h00;
    ff_ram[15201] = 8'h00;
    ff_ram[15202] = 8'h00;
    ff_ram[15203] = 8'h00;
    ff_ram[15204] = 8'h00;
    ff_ram[15205] = 8'h00;
    ff_ram[15206] = 8'h00;
    ff_ram[15207] = 8'h00;
    ff_ram[15208] = 8'h00;
    ff_ram[15209] = 8'h00;
    ff_ram[15210] = 8'h00;
    ff_ram[15211] = 8'h00;
    ff_ram[15212] = 8'h00;
    ff_ram[15213] = 8'h00;
    ff_ram[15214] = 8'h00;
    ff_ram[15215] = 8'h00;
    ff_ram[15216] = 8'h00;
    ff_ram[15217] = 8'h00;
    ff_ram[15218] = 8'h00;
    ff_ram[15219] = 8'h00;
    ff_ram[15220] = 8'h00;
    ff_ram[15221] = 8'h00;
    ff_ram[15222] = 8'h00;
    ff_ram[15223] = 8'h00;
    ff_ram[15224] = 8'h00;
    ff_ram[15225] = 8'h00;
    ff_ram[15226] = 8'h00;
    ff_ram[15227] = 8'h00;
    ff_ram[15228] = 8'h00;
    ff_ram[15229] = 8'h00;
    ff_ram[15230] = 8'h00;
    ff_ram[15231] = 8'h00;
    ff_ram[15232] = 8'h00;
    ff_ram[15233] = 8'h00;
    ff_ram[15234] = 8'h00;
    ff_ram[15235] = 8'h00;
    ff_ram[15236] = 8'h00;
    ff_ram[15237] = 8'h00;
    ff_ram[15238] = 8'h00;
    ff_ram[15239] = 8'h00;
    ff_ram[15240] = 8'h00;
    ff_ram[15241] = 8'h00;
    ff_ram[15242] = 8'h00;
    ff_ram[15243] = 8'h00;
    ff_ram[15244] = 8'h00;
    ff_ram[15245] = 8'h00;
    ff_ram[15246] = 8'h00;
    ff_ram[15247] = 8'h00;
    ff_ram[15248] = 8'h00;
    ff_ram[15249] = 8'h00;
    ff_ram[15250] = 8'h00;
    ff_ram[15251] = 8'h00;
    ff_ram[15252] = 8'h00;
    ff_ram[15253] = 8'h00;
    ff_ram[15254] = 8'h00;
    ff_ram[15255] = 8'h00;
    ff_ram[15256] = 8'h00;
    ff_ram[15257] = 8'h00;
    ff_ram[15258] = 8'h00;
    ff_ram[15259] = 8'h00;
    ff_ram[15260] = 8'h00;
    ff_ram[15261] = 8'h00;
    ff_ram[15262] = 8'h00;
    ff_ram[15263] = 8'h00;
    ff_ram[15264] = 8'h00;
    ff_ram[15265] = 8'h00;
    ff_ram[15266] = 8'h00;
    ff_ram[15267] = 8'h00;
    ff_ram[15268] = 8'h00;
    ff_ram[15269] = 8'h00;
    ff_ram[15270] = 8'h00;
    ff_ram[15271] = 8'h00;
    ff_ram[15272] = 8'h00;
    ff_ram[15273] = 8'h00;
    ff_ram[15274] = 8'h00;
    ff_ram[15275] = 8'h00;
    ff_ram[15276] = 8'h00;
    ff_ram[15277] = 8'h00;
    ff_ram[15278] = 8'h00;
    ff_ram[15279] = 8'h00;
    ff_ram[15280] = 8'h00;
    ff_ram[15281] = 8'h00;
    ff_ram[15282] = 8'h00;
    ff_ram[15283] = 8'h00;
    ff_ram[15284] = 8'h00;
    ff_ram[15285] = 8'h00;
    ff_ram[15286] = 8'h00;
    ff_ram[15287] = 8'h00;
    ff_ram[15288] = 8'h00;
    ff_ram[15289] = 8'h00;
    ff_ram[15290] = 8'h00;
    ff_ram[15291] = 8'h00;
    ff_ram[15292] = 8'h00;
    ff_ram[15293] = 8'h00;
    ff_ram[15294] = 8'h00;
    ff_ram[15295] = 8'h00;
    ff_ram[15296] = 8'h00;
    ff_ram[15297] = 8'h00;
    ff_ram[15298] = 8'h00;
    ff_ram[15299] = 8'h00;
    ff_ram[15300] = 8'h00;
    ff_ram[15301] = 8'h00;
    ff_ram[15302] = 8'h00;
    ff_ram[15303] = 8'h00;
    ff_ram[15304] = 8'h00;
    ff_ram[15305] = 8'h00;
    ff_ram[15306] = 8'h00;
    ff_ram[15307] = 8'h00;
    ff_ram[15308] = 8'h00;
    ff_ram[15309] = 8'h00;
    ff_ram[15310] = 8'h00;
    ff_ram[15311] = 8'h00;
    ff_ram[15312] = 8'h00;
    ff_ram[15313] = 8'h00;
    ff_ram[15314] = 8'h00;
    ff_ram[15315] = 8'h00;
    ff_ram[15316] = 8'h00;
    ff_ram[15317] = 8'h00;
    ff_ram[15318] = 8'h00;
    ff_ram[15319] = 8'h00;
    ff_ram[15320] = 8'h00;
    ff_ram[15321] = 8'h00;
    ff_ram[15322] = 8'h00;
    ff_ram[15323] = 8'h00;
    ff_ram[15324] = 8'h00;
    ff_ram[15325] = 8'h00;
    ff_ram[15326] = 8'h00;
    ff_ram[15327] = 8'h00;
    ff_ram[15328] = 8'h00;
    ff_ram[15329] = 8'h00;
    ff_ram[15330] = 8'h00;
    ff_ram[15331] = 8'h00;
    ff_ram[15332] = 8'h00;
    ff_ram[15333] = 8'h00;
    ff_ram[15334] = 8'h00;
    ff_ram[15335] = 8'h00;
    ff_ram[15336] = 8'h00;
    ff_ram[15337] = 8'h00;
    ff_ram[15338] = 8'h00;
    ff_ram[15339] = 8'h00;
    ff_ram[15340] = 8'h00;
    ff_ram[15341] = 8'h00;
    ff_ram[15342] = 8'h00;
    ff_ram[15343] = 8'h00;
    ff_ram[15344] = 8'h00;
    ff_ram[15345] = 8'h00;
    ff_ram[15346] = 8'h00;
    ff_ram[15347] = 8'h00;
    ff_ram[15348] = 8'h00;
    ff_ram[15349] = 8'h00;
    ff_ram[15350] = 8'h00;
    ff_ram[15351] = 8'h00;
    ff_ram[15352] = 8'h00;
    ff_ram[15353] = 8'h00;
    ff_ram[15354] = 8'h00;
    ff_ram[15355] = 8'h00;
    ff_ram[15356] = 8'h00;
    ff_ram[15357] = 8'h00;
    ff_ram[15358] = 8'h00;
    ff_ram[15359] = 8'h00;
    ff_ram[15360] = 8'h00;
    ff_ram[15361] = 8'h00;
    ff_ram[15362] = 8'h00;
    ff_ram[15363] = 8'h00;
    ff_ram[15364] = 8'h00;
    ff_ram[15365] = 8'h00;
    ff_ram[15366] = 8'h00;
    ff_ram[15367] = 8'h00;
    ff_ram[15368] = 8'h00;
    ff_ram[15369] = 8'h00;
    ff_ram[15370] = 8'h00;
    ff_ram[15371] = 8'h00;
    ff_ram[15372] = 8'h00;
    ff_ram[15373] = 8'h00;
    ff_ram[15374] = 8'h00;
    ff_ram[15375] = 8'h00;
    ff_ram[15376] = 8'h00;
    ff_ram[15377] = 8'h00;
    ff_ram[15378] = 8'h00;
    ff_ram[15379] = 8'h00;
    ff_ram[15380] = 8'h00;
    ff_ram[15381] = 8'h00;
    ff_ram[15382] = 8'h00;
    ff_ram[15383] = 8'h00;
    ff_ram[15384] = 8'h00;
    ff_ram[15385] = 8'h00;
    ff_ram[15386] = 8'h00;
    ff_ram[15387] = 8'h00;
    ff_ram[15388] = 8'h00;
    ff_ram[15389] = 8'h00;
    ff_ram[15390] = 8'h00;
    ff_ram[15391] = 8'h00;
    ff_ram[15392] = 8'h00;
    ff_ram[15393] = 8'h00;
    ff_ram[15394] = 8'h00;
    ff_ram[15395] = 8'h00;
    ff_ram[15396] = 8'h00;
    ff_ram[15397] = 8'h00;
    ff_ram[15398] = 8'h00;
    ff_ram[15399] = 8'h00;
    ff_ram[15400] = 8'h00;
    ff_ram[15401] = 8'h00;
    ff_ram[15402] = 8'h00;
    ff_ram[15403] = 8'h00;
    ff_ram[15404] = 8'h00;
    ff_ram[15405] = 8'h00;
    ff_ram[15406] = 8'h00;
    ff_ram[15407] = 8'h00;
    ff_ram[15408] = 8'h00;
    ff_ram[15409] = 8'h00;
    ff_ram[15410] = 8'h00;
    ff_ram[15411] = 8'h00;
    ff_ram[15412] = 8'h00;
    ff_ram[15413] = 8'h00;
    ff_ram[15414] = 8'h00;
    ff_ram[15415] = 8'h00;
    ff_ram[15416] = 8'h00;
    ff_ram[15417] = 8'h00;
    ff_ram[15418] = 8'h00;
    ff_ram[15419] = 8'h00;
    ff_ram[15420] = 8'h00;
    ff_ram[15421] = 8'h00;
    ff_ram[15422] = 8'h00;
    ff_ram[15423] = 8'h00;
    ff_ram[15424] = 8'h00;
    ff_ram[15425] = 8'h00;
    ff_ram[15426] = 8'h00;
    ff_ram[15427] = 8'h00;
    ff_ram[15428] = 8'h00;
    ff_ram[15429] = 8'h00;
    ff_ram[15430] = 8'h00;
    ff_ram[15431] = 8'h00;
    ff_ram[15432] = 8'h00;
    ff_ram[15433] = 8'h00;
    ff_ram[15434] = 8'h00;
    ff_ram[15435] = 8'h00;
    ff_ram[15436] = 8'h00;
    ff_ram[15437] = 8'h00;
    ff_ram[15438] = 8'h00;
    ff_ram[15439] = 8'h00;
    ff_ram[15440] = 8'h00;
    ff_ram[15441] = 8'h00;
    ff_ram[15442] = 8'h00;
    ff_ram[15443] = 8'h00;
    ff_ram[15444] = 8'h00;
    ff_ram[15445] = 8'h00;
    ff_ram[15446] = 8'h00;
    ff_ram[15447] = 8'h00;
    ff_ram[15448] = 8'h00;
    ff_ram[15449] = 8'h00;
    ff_ram[15450] = 8'h00;
    ff_ram[15451] = 8'h00;
    ff_ram[15452] = 8'h00;
    ff_ram[15453] = 8'h00;
    ff_ram[15454] = 8'h00;
    ff_ram[15455] = 8'h00;
    ff_ram[15456] = 8'h00;
    ff_ram[15457] = 8'h00;
    ff_ram[15458] = 8'h00;
    ff_ram[15459] = 8'h00;
    ff_ram[15460] = 8'h00;
    ff_ram[15461] = 8'h00;
    ff_ram[15462] = 8'h00;
    ff_ram[15463] = 8'h00;
    ff_ram[15464] = 8'h00;
    ff_ram[15465] = 8'h00;
    ff_ram[15466] = 8'h00;
    ff_ram[15467] = 8'h00;
    ff_ram[15468] = 8'h00;
    ff_ram[15469] = 8'h00;
    ff_ram[15470] = 8'h00;
    ff_ram[15471] = 8'h00;
    ff_ram[15472] = 8'h00;
    ff_ram[15473] = 8'h00;
    ff_ram[15474] = 8'h00;
    ff_ram[15475] = 8'h00;
    ff_ram[15476] = 8'h00;
    ff_ram[15477] = 8'h00;
    ff_ram[15478] = 8'h00;
    ff_ram[15479] = 8'h00;
    ff_ram[15480] = 8'h00;
    ff_ram[15481] = 8'h00;
    ff_ram[15482] = 8'h00;
    ff_ram[15483] = 8'h00;
    ff_ram[15484] = 8'h00;
    ff_ram[15485] = 8'h00;
    ff_ram[15486] = 8'h00;
    ff_ram[15487] = 8'h00;
    ff_ram[15488] = 8'h00;
    ff_ram[15489] = 8'h00;
    ff_ram[15490] = 8'h00;
    ff_ram[15491] = 8'h00;
    ff_ram[15492] = 8'h00;
    ff_ram[15493] = 8'h00;
    ff_ram[15494] = 8'h00;
    ff_ram[15495] = 8'h00;
    ff_ram[15496] = 8'h00;
    ff_ram[15497] = 8'h00;
    ff_ram[15498] = 8'h00;
    ff_ram[15499] = 8'h00;
    ff_ram[15500] = 8'h00;
    ff_ram[15501] = 8'h00;
    ff_ram[15502] = 8'h00;
    ff_ram[15503] = 8'h00;
    ff_ram[15504] = 8'h00;
    ff_ram[15505] = 8'h00;
    ff_ram[15506] = 8'h00;
    ff_ram[15507] = 8'h00;
    ff_ram[15508] = 8'h00;
    ff_ram[15509] = 8'h00;
    ff_ram[15510] = 8'h00;
    ff_ram[15511] = 8'h00;
    ff_ram[15512] = 8'h00;
    ff_ram[15513] = 8'h00;
    ff_ram[15514] = 8'h00;
    ff_ram[15515] = 8'h00;
    ff_ram[15516] = 8'h00;
    ff_ram[15517] = 8'h00;
    ff_ram[15518] = 8'h00;
    ff_ram[15519] = 8'h00;
    ff_ram[15520] = 8'h00;
    ff_ram[15521] = 8'h00;
    ff_ram[15522] = 8'h00;
    ff_ram[15523] = 8'h00;
    ff_ram[15524] = 8'h00;
    ff_ram[15525] = 8'h00;
    ff_ram[15526] = 8'h00;
    ff_ram[15527] = 8'h00;
    ff_ram[15528] = 8'h00;
    ff_ram[15529] = 8'h00;
    ff_ram[15530] = 8'h00;
    ff_ram[15531] = 8'h00;
    ff_ram[15532] = 8'h00;
    ff_ram[15533] = 8'h00;
    ff_ram[15534] = 8'h00;
    ff_ram[15535] = 8'h00;
    ff_ram[15536] = 8'h00;
    ff_ram[15537] = 8'h00;
    ff_ram[15538] = 8'h00;
    ff_ram[15539] = 8'h00;
    ff_ram[15540] = 8'h00;
    ff_ram[15541] = 8'h00;
    ff_ram[15542] = 8'h00;
    ff_ram[15543] = 8'h00;
    ff_ram[15544] = 8'h00;
    ff_ram[15545] = 8'h00;
    ff_ram[15546] = 8'h00;
    ff_ram[15547] = 8'h00;
    ff_ram[15548] = 8'h00;
    ff_ram[15549] = 8'h00;
    ff_ram[15550] = 8'h00;
    ff_ram[15551] = 8'h00;
    ff_ram[15552] = 8'h00;
    ff_ram[15553] = 8'h00;
    ff_ram[15554] = 8'h00;
    ff_ram[15555] = 8'h00;
    ff_ram[15556] = 8'h00;
    ff_ram[15557] = 8'h00;
    ff_ram[15558] = 8'h00;
    ff_ram[15559] = 8'h00;
    ff_ram[15560] = 8'h00;
    ff_ram[15561] = 8'h00;
    ff_ram[15562] = 8'h00;
    ff_ram[15563] = 8'h00;
    ff_ram[15564] = 8'h00;
    ff_ram[15565] = 8'h00;
    ff_ram[15566] = 8'h00;
    ff_ram[15567] = 8'h00;
    ff_ram[15568] = 8'h00;
    ff_ram[15569] = 8'h00;
    ff_ram[15570] = 8'h00;
    ff_ram[15571] = 8'h00;
    ff_ram[15572] = 8'h00;
    ff_ram[15573] = 8'h00;
    ff_ram[15574] = 8'h00;
    ff_ram[15575] = 8'h00;
    ff_ram[15576] = 8'h00;
    ff_ram[15577] = 8'h00;
    ff_ram[15578] = 8'h00;
    ff_ram[15579] = 8'h00;
    ff_ram[15580] = 8'h00;
    ff_ram[15581] = 8'h00;
    ff_ram[15582] = 8'h00;
    ff_ram[15583] = 8'h00;
    ff_ram[15584] = 8'h00;
    ff_ram[15585] = 8'h00;
    ff_ram[15586] = 8'h00;
    ff_ram[15587] = 8'h00;
    ff_ram[15588] = 8'h00;
    ff_ram[15589] = 8'h00;
    ff_ram[15590] = 8'h00;
    ff_ram[15591] = 8'h00;
    ff_ram[15592] = 8'h00;
    ff_ram[15593] = 8'h00;
    ff_ram[15594] = 8'h00;
    ff_ram[15595] = 8'h00;
    ff_ram[15596] = 8'h00;
    ff_ram[15597] = 8'h00;
    ff_ram[15598] = 8'h00;
    ff_ram[15599] = 8'h00;
    ff_ram[15600] = 8'h00;
    ff_ram[15601] = 8'h00;
    ff_ram[15602] = 8'h00;
    ff_ram[15603] = 8'h00;
    ff_ram[15604] = 8'h00;
    ff_ram[15605] = 8'h00;
    ff_ram[15606] = 8'h00;
    ff_ram[15607] = 8'h00;
    ff_ram[15608] = 8'h00;
    ff_ram[15609] = 8'h00;
    ff_ram[15610] = 8'h00;
    ff_ram[15611] = 8'h00;
    ff_ram[15612] = 8'h00;
    ff_ram[15613] = 8'h00;
    ff_ram[15614] = 8'h00;
    ff_ram[15615] = 8'h00;
    ff_ram[15616] = 8'h00;
    ff_ram[15617] = 8'h00;
    ff_ram[15618] = 8'h00;
    ff_ram[15619] = 8'h00;
    ff_ram[15620] = 8'h00;
    ff_ram[15621] = 8'h00;
    ff_ram[15622] = 8'h00;
    ff_ram[15623] = 8'h00;
    ff_ram[15624] = 8'h00;
    ff_ram[15625] = 8'h00;
    ff_ram[15626] = 8'h00;
    ff_ram[15627] = 8'h00;
    ff_ram[15628] = 8'h00;
    ff_ram[15629] = 8'h00;
    ff_ram[15630] = 8'h00;
    ff_ram[15631] = 8'h00;
    ff_ram[15632] = 8'h00;
    ff_ram[15633] = 8'h00;
    ff_ram[15634] = 8'h00;
    ff_ram[15635] = 8'h00;
    ff_ram[15636] = 8'h00;
    ff_ram[15637] = 8'h00;
    ff_ram[15638] = 8'h00;
    ff_ram[15639] = 8'h00;
    ff_ram[15640] = 8'h00;
    ff_ram[15641] = 8'h00;
    ff_ram[15642] = 8'h00;
    ff_ram[15643] = 8'h00;
    ff_ram[15644] = 8'h00;
    ff_ram[15645] = 8'h00;
    ff_ram[15646] = 8'h00;
    ff_ram[15647] = 8'h00;
    ff_ram[15648] = 8'h00;
    ff_ram[15649] = 8'h00;
    ff_ram[15650] = 8'h00;
    ff_ram[15651] = 8'h00;
    ff_ram[15652] = 8'h00;
    ff_ram[15653] = 8'h00;
    ff_ram[15654] = 8'h00;
    ff_ram[15655] = 8'h00;
    ff_ram[15656] = 8'h00;
    ff_ram[15657] = 8'h00;
    ff_ram[15658] = 8'h00;
    ff_ram[15659] = 8'h00;
    ff_ram[15660] = 8'h00;
    ff_ram[15661] = 8'h00;
    ff_ram[15662] = 8'h00;
    ff_ram[15663] = 8'h00;
    ff_ram[15664] = 8'h00;
    ff_ram[15665] = 8'h00;
    ff_ram[15666] = 8'h00;
    ff_ram[15667] = 8'h00;
    ff_ram[15668] = 8'h00;
    ff_ram[15669] = 8'h00;
    ff_ram[15670] = 8'h00;
    ff_ram[15671] = 8'h00;
    ff_ram[15672] = 8'h00;
    ff_ram[15673] = 8'h00;
    ff_ram[15674] = 8'h00;
    ff_ram[15675] = 8'h00;
    ff_ram[15676] = 8'h00;
    ff_ram[15677] = 8'h00;
    ff_ram[15678] = 8'h00;
    ff_ram[15679] = 8'h00;
    ff_ram[15680] = 8'h00;
    ff_ram[15681] = 8'h00;
    ff_ram[15682] = 8'h00;
    ff_ram[15683] = 8'h00;
    ff_ram[15684] = 8'h00;
    ff_ram[15685] = 8'h00;
    ff_ram[15686] = 8'h00;
    ff_ram[15687] = 8'h00;
    ff_ram[15688] = 8'h00;
    ff_ram[15689] = 8'h00;
    ff_ram[15690] = 8'h00;
    ff_ram[15691] = 8'h00;
    ff_ram[15692] = 8'h00;
    ff_ram[15693] = 8'h00;
    ff_ram[15694] = 8'h00;
    ff_ram[15695] = 8'h00;
    ff_ram[15696] = 8'h00;
    ff_ram[15697] = 8'h00;
    ff_ram[15698] = 8'h00;
    ff_ram[15699] = 8'h00;
    ff_ram[15700] = 8'h00;
    ff_ram[15701] = 8'h00;
    ff_ram[15702] = 8'h00;
    ff_ram[15703] = 8'h00;
    ff_ram[15704] = 8'h00;
    ff_ram[15705] = 8'h00;
    ff_ram[15706] = 8'h00;
    ff_ram[15707] = 8'h00;
    ff_ram[15708] = 8'h00;
    ff_ram[15709] = 8'h00;
    ff_ram[15710] = 8'h00;
    ff_ram[15711] = 8'h00;
    ff_ram[15712] = 8'h00;
    ff_ram[15713] = 8'h00;
    ff_ram[15714] = 8'h00;
    ff_ram[15715] = 8'h00;
    ff_ram[15716] = 8'h00;
    ff_ram[15717] = 8'h00;
    ff_ram[15718] = 8'h00;
    ff_ram[15719] = 8'h00;
    ff_ram[15720] = 8'h00;
    ff_ram[15721] = 8'h00;
    ff_ram[15722] = 8'h00;
    ff_ram[15723] = 8'h00;
    ff_ram[15724] = 8'h00;
    ff_ram[15725] = 8'h00;
    ff_ram[15726] = 8'h00;
    ff_ram[15727] = 8'h00;
    ff_ram[15728] = 8'h00;
    ff_ram[15729] = 8'h00;
    ff_ram[15730] = 8'h00;
    ff_ram[15731] = 8'h00;
    ff_ram[15732] = 8'h00;
    ff_ram[15733] = 8'h00;
    ff_ram[15734] = 8'h00;
    ff_ram[15735] = 8'h00;
    ff_ram[15736] = 8'h00;
    ff_ram[15737] = 8'h00;
    ff_ram[15738] = 8'h00;
    ff_ram[15739] = 8'h00;
    ff_ram[15740] = 8'h00;
    ff_ram[15741] = 8'h00;
    ff_ram[15742] = 8'h00;
    ff_ram[15743] = 8'h00;
    ff_ram[15744] = 8'h00;
    ff_ram[15745] = 8'h00;
    ff_ram[15746] = 8'h00;
    ff_ram[15747] = 8'h00;
    ff_ram[15748] = 8'h00;
    ff_ram[15749] = 8'h00;
    ff_ram[15750] = 8'h00;
    ff_ram[15751] = 8'h00;
    ff_ram[15752] = 8'h00;
    ff_ram[15753] = 8'h00;
    ff_ram[15754] = 8'h00;
    ff_ram[15755] = 8'h00;
    ff_ram[15756] = 8'h00;
    ff_ram[15757] = 8'h00;
    ff_ram[15758] = 8'h00;
    ff_ram[15759] = 8'h00;
    ff_ram[15760] = 8'h00;
    ff_ram[15761] = 8'h00;
    ff_ram[15762] = 8'h00;
    ff_ram[15763] = 8'h00;
    ff_ram[15764] = 8'h00;
    ff_ram[15765] = 8'h00;
    ff_ram[15766] = 8'h00;
    ff_ram[15767] = 8'h00;
    ff_ram[15768] = 8'h00;
    ff_ram[15769] = 8'h00;
    ff_ram[15770] = 8'h00;
    ff_ram[15771] = 8'h00;
    ff_ram[15772] = 8'h00;
    ff_ram[15773] = 8'h00;
    ff_ram[15774] = 8'h00;
    ff_ram[15775] = 8'h00;
    ff_ram[15776] = 8'h00;
    ff_ram[15777] = 8'h00;
    ff_ram[15778] = 8'h00;
    ff_ram[15779] = 8'h00;
    ff_ram[15780] = 8'h00;
    ff_ram[15781] = 8'h00;
    ff_ram[15782] = 8'h00;
    ff_ram[15783] = 8'h00;
    ff_ram[15784] = 8'h00;
    ff_ram[15785] = 8'h00;
    ff_ram[15786] = 8'h00;
    ff_ram[15787] = 8'h00;
    ff_ram[15788] = 8'h00;
    ff_ram[15789] = 8'h00;
    ff_ram[15790] = 8'h00;
    ff_ram[15791] = 8'h00;
    ff_ram[15792] = 8'h00;
    ff_ram[15793] = 8'h00;
    ff_ram[15794] = 8'h00;
    ff_ram[15795] = 8'h00;
    ff_ram[15796] = 8'h00;
    ff_ram[15797] = 8'h00;
    ff_ram[15798] = 8'h00;
    ff_ram[15799] = 8'h00;
    ff_ram[15800] = 8'h00;
    ff_ram[15801] = 8'h00;
    ff_ram[15802] = 8'h00;
    ff_ram[15803] = 8'h00;
    ff_ram[15804] = 8'h00;
    ff_ram[15805] = 8'h00;
    ff_ram[15806] = 8'h00;
    ff_ram[15807] = 8'h00;
    ff_ram[15808] = 8'h00;
    ff_ram[15809] = 8'h00;
    ff_ram[15810] = 8'h00;
    ff_ram[15811] = 8'h00;
    ff_ram[15812] = 8'h00;
    ff_ram[15813] = 8'h00;
    ff_ram[15814] = 8'h00;
    ff_ram[15815] = 8'h00;
    ff_ram[15816] = 8'h00;
    ff_ram[15817] = 8'h00;
    ff_ram[15818] = 8'h00;
    ff_ram[15819] = 8'h00;
    ff_ram[15820] = 8'h00;
    ff_ram[15821] = 8'h00;
    ff_ram[15822] = 8'h00;
    ff_ram[15823] = 8'h00;
    ff_ram[15824] = 8'h00;
    ff_ram[15825] = 8'h00;
    ff_ram[15826] = 8'h00;
    ff_ram[15827] = 8'h00;
    ff_ram[15828] = 8'h00;
    ff_ram[15829] = 8'h00;
    ff_ram[15830] = 8'h00;
    ff_ram[15831] = 8'h00;
    ff_ram[15832] = 8'h00;
    ff_ram[15833] = 8'h00;
    ff_ram[15834] = 8'h00;
    ff_ram[15835] = 8'h00;
    ff_ram[15836] = 8'h00;
    ff_ram[15837] = 8'h00;
    ff_ram[15838] = 8'h00;
    ff_ram[15839] = 8'h00;
    ff_ram[15840] = 8'h00;
    ff_ram[15841] = 8'h00;
    ff_ram[15842] = 8'h00;
    ff_ram[15843] = 8'h00;
    ff_ram[15844] = 8'h00;
    ff_ram[15845] = 8'h00;
    ff_ram[15846] = 8'h00;
    ff_ram[15847] = 8'h00;
    ff_ram[15848] = 8'h00;
    ff_ram[15849] = 8'h00;
    ff_ram[15850] = 8'h00;
    ff_ram[15851] = 8'h00;
    ff_ram[15852] = 8'h00;
    ff_ram[15853] = 8'h00;
    ff_ram[15854] = 8'h00;
    ff_ram[15855] = 8'h00;
    ff_ram[15856] = 8'h00;
    ff_ram[15857] = 8'h00;
    ff_ram[15858] = 8'h00;
    ff_ram[15859] = 8'h00;
    ff_ram[15860] = 8'h00;
    ff_ram[15861] = 8'h00;
    ff_ram[15862] = 8'h00;
    ff_ram[15863] = 8'h00;
    ff_ram[15864] = 8'h00;
    ff_ram[15865] = 8'h00;
    ff_ram[15866] = 8'h00;
    ff_ram[15867] = 8'h00;
    ff_ram[15868] = 8'h00;
    ff_ram[15869] = 8'h00;
    ff_ram[15870] = 8'h00;
    ff_ram[15871] = 8'h00;
    ff_ram[15872] = 8'h00;
    ff_ram[15873] = 8'h00;
    ff_ram[15874] = 8'h00;
    ff_ram[15875] = 8'h00;
    ff_ram[15876] = 8'h00;
    ff_ram[15877] = 8'h00;
    ff_ram[15878] = 8'h00;
    ff_ram[15879] = 8'h00;
    ff_ram[15880] = 8'h00;
    ff_ram[15881] = 8'h00;
    ff_ram[15882] = 8'h00;
    ff_ram[15883] = 8'h00;
    ff_ram[15884] = 8'h00;
    ff_ram[15885] = 8'h00;
    ff_ram[15886] = 8'h00;
    ff_ram[15887] = 8'h00;
    ff_ram[15888] = 8'h00;
    ff_ram[15889] = 8'h00;
    ff_ram[15890] = 8'h00;
    ff_ram[15891] = 8'h00;
    ff_ram[15892] = 8'h00;
    ff_ram[15893] = 8'h00;
    ff_ram[15894] = 8'h00;
    ff_ram[15895] = 8'h00;
    ff_ram[15896] = 8'h00;
    ff_ram[15897] = 8'h00;
    ff_ram[15898] = 8'h00;
    ff_ram[15899] = 8'h00;
    ff_ram[15900] = 8'h00;
    ff_ram[15901] = 8'h00;
    ff_ram[15902] = 8'h00;
    ff_ram[15903] = 8'h00;
    ff_ram[15904] = 8'h00;
    ff_ram[15905] = 8'h00;
    ff_ram[15906] = 8'h00;
    ff_ram[15907] = 8'h00;
    ff_ram[15908] = 8'h00;
    ff_ram[15909] = 8'h00;
    ff_ram[15910] = 8'h00;
    ff_ram[15911] = 8'h00;
    ff_ram[15912] = 8'h00;
    ff_ram[15913] = 8'h00;
    ff_ram[15914] = 8'h00;
    ff_ram[15915] = 8'h00;
    ff_ram[15916] = 8'h00;
    ff_ram[15917] = 8'h00;
    ff_ram[15918] = 8'h00;
    ff_ram[15919] = 8'h00;
    ff_ram[15920] = 8'h00;
    ff_ram[15921] = 8'h00;
    ff_ram[15922] = 8'h00;
    ff_ram[15923] = 8'h00;
    ff_ram[15924] = 8'h00;
    ff_ram[15925] = 8'h00;
    ff_ram[15926] = 8'h00;
    ff_ram[15927] = 8'h00;
    ff_ram[15928] = 8'h00;
    ff_ram[15929] = 8'h00;
    ff_ram[15930] = 8'h00;
    ff_ram[15931] = 8'h00;
    ff_ram[15932] = 8'h00;
    ff_ram[15933] = 8'h00;
    ff_ram[15934] = 8'h00;
    ff_ram[15935] = 8'h00;
    ff_ram[15936] = 8'h00;
    ff_ram[15937] = 8'h00;
    ff_ram[15938] = 8'h00;
    ff_ram[15939] = 8'h00;
    ff_ram[15940] = 8'h00;
    ff_ram[15941] = 8'h00;
    ff_ram[15942] = 8'h00;
    ff_ram[15943] = 8'h00;
    ff_ram[15944] = 8'h00;
    ff_ram[15945] = 8'h00;
    ff_ram[15946] = 8'h00;
    ff_ram[15947] = 8'h00;
    ff_ram[15948] = 8'h00;
    ff_ram[15949] = 8'h00;
    ff_ram[15950] = 8'h00;
    ff_ram[15951] = 8'h00;
    ff_ram[15952] = 8'h00;
    ff_ram[15953] = 8'h00;
    ff_ram[15954] = 8'h00;
    ff_ram[15955] = 8'h00;
    ff_ram[15956] = 8'h00;
    ff_ram[15957] = 8'h00;
    ff_ram[15958] = 8'h00;
    ff_ram[15959] = 8'h00;
    ff_ram[15960] = 8'h00;
    ff_ram[15961] = 8'h00;
    ff_ram[15962] = 8'h00;
    ff_ram[15963] = 8'h00;
    ff_ram[15964] = 8'h00;
    ff_ram[15965] = 8'h00;
    ff_ram[15966] = 8'h00;
    ff_ram[15967] = 8'h00;
    ff_ram[15968] = 8'h00;
    ff_ram[15969] = 8'h00;
    ff_ram[15970] = 8'h00;
    ff_ram[15971] = 8'h00;
    ff_ram[15972] = 8'h00;
    ff_ram[15973] = 8'h00;
    ff_ram[15974] = 8'h00;
    ff_ram[15975] = 8'h00;
    ff_ram[15976] = 8'h00;
    ff_ram[15977] = 8'h00;
    ff_ram[15978] = 8'h00;
    ff_ram[15979] = 8'h00;
    ff_ram[15980] = 8'h00;
    ff_ram[15981] = 8'h00;
    ff_ram[15982] = 8'h00;
    ff_ram[15983] = 8'h00;
    ff_ram[15984] = 8'h00;
    ff_ram[15985] = 8'h00;
    ff_ram[15986] = 8'h00;
    ff_ram[15987] = 8'h00;
    ff_ram[15988] = 8'h00;
    ff_ram[15989] = 8'h00;
    ff_ram[15990] = 8'h00;
    ff_ram[15991] = 8'h00;
    ff_ram[15992] = 8'h00;
    ff_ram[15993] = 8'h00;
    ff_ram[15994] = 8'h00;
    ff_ram[15995] = 8'h00;
    ff_ram[15996] = 8'h00;
    ff_ram[15997] = 8'h00;
    ff_ram[15998] = 8'h00;
    ff_ram[15999] = 8'h00;
    ff_ram[16000] = 8'h00;
    ff_ram[16001] = 8'h00;
    ff_ram[16002] = 8'h00;
    ff_ram[16003] = 8'h00;
    ff_ram[16004] = 8'h00;
    ff_ram[16005] = 8'h00;
    ff_ram[16006] = 8'h00;
    ff_ram[16007] = 8'h00;
    ff_ram[16008] = 8'h00;
    ff_ram[16009] = 8'h00;
    ff_ram[16010] = 8'h00;
    ff_ram[16011] = 8'h00;
    ff_ram[16012] = 8'h00;
    ff_ram[16013] = 8'h00;
    ff_ram[16014] = 8'h00;
    ff_ram[16015] = 8'h00;
    ff_ram[16016] = 8'h00;
    ff_ram[16017] = 8'h00;
    ff_ram[16018] = 8'h00;
    ff_ram[16019] = 8'h00;
    ff_ram[16020] = 8'h00;
    ff_ram[16021] = 8'h00;
    ff_ram[16022] = 8'h00;
    ff_ram[16023] = 8'h00;
    ff_ram[16024] = 8'h00;
    ff_ram[16025] = 8'h00;
    ff_ram[16026] = 8'h00;
    ff_ram[16027] = 8'h00;
    ff_ram[16028] = 8'h00;
    ff_ram[16029] = 8'h00;
    ff_ram[16030] = 8'h00;
    ff_ram[16031] = 8'h00;
    ff_ram[16032] = 8'h00;
    ff_ram[16033] = 8'h00;
    ff_ram[16034] = 8'h00;
    ff_ram[16035] = 8'h00;
    ff_ram[16036] = 8'h00;
    ff_ram[16037] = 8'h00;
    ff_ram[16038] = 8'h00;
    ff_ram[16039] = 8'h00;
    ff_ram[16040] = 8'h00;
    ff_ram[16041] = 8'h00;
    ff_ram[16042] = 8'h00;
    ff_ram[16043] = 8'h00;
    ff_ram[16044] = 8'h00;
    ff_ram[16045] = 8'h00;
    ff_ram[16046] = 8'h00;
    ff_ram[16047] = 8'h00;
    ff_ram[16048] = 8'h00;
    ff_ram[16049] = 8'h00;
    ff_ram[16050] = 8'h00;
    ff_ram[16051] = 8'h00;
    ff_ram[16052] = 8'h00;
    ff_ram[16053] = 8'h00;
    ff_ram[16054] = 8'h00;
    ff_ram[16055] = 8'h00;
    ff_ram[16056] = 8'h00;
    ff_ram[16057] = 8'h00;
    ff_ram[16058] = 8'h00;
    ff_ram[16059] = 8'h00;
    ff_ram[16060] = 8'h00;
    ff_ram[16061] = 8'h00;
    ff_ram[16062] = 8'h00;
    ff_ram[16063] = 8'h00;
    ff_ram[16064] = 8'h00;
    ff_ram[16065] = 8'h00;
    ff_ram[16066] = 8'h00;
    ff_ram[16067] = 8'h00;
    ff_ram[16068] = 8'h00;
    ff_ram[16069] = 8'h00;
    ff_ram[16070] = 8'h00;
    ff_ram[16071] = 8'h00;
    ff_ram[16072] = 8'h00;
    ff_ram[16073] = 8'h00;
    ff_ram[16074] = 8'h00;
    ff_ram[16075] = 8'h00;
    ff_ram[16076] = 8'h00;
    ff_ram[16077] = 8'h00;
    ff_ram[16078] = 8'h00;
    ff_ram[16079] = 8'h00;
    ff_ram[16080] = 8'h00;
    ff_ram[16081] = 8'h00;
    ff_ram[16082] = 8'h00;
    ff_ram[16083] = 8'h00;
    ff_ram[16084] = 8'h00;
    ff_ram[16085] = 8'h00;
    ff_ram[16086] = 8'h00;
    ff_ram[16087] = 8'h00;
    ff_ram[16088] = 8'h00;
    ff_ram[16089] = 8'h00;
    ff_ram[16090] = 8'h00;
    ff_ram[16091] = 8'h00;
    ff_ram[16092] = 8'h00;
    ff_ram[16093] = 8'h00;
    ff_ram[16094] = 8'h00;
    ff_ram[16095] = 8'h00;
    ff_ram[16096] = 8'h00;
    ff_ram[16097] = 8'h00;
    ff_ram[16098] = 8'h00;
    ff_ram[16099] = 8'h00;
    ff_ram[16100] = 8'h00;
    ff_ram[16101] = 8'h00;
    ff_ram[16102] = 8'h00;
    ff_ram[16103] = 8'h00;
    ff_ram[16104] = 8'h00;
    ff_ram[16105] = 8'h00;
    ff_ram[16106] = 8'h00;
    ff_ram[16107] = 8'h00;
    ff_ram[16108] = 8'h00;
    ff_ram[16109] = 8'h00;
    ff_ram[16110] = 8'h00;
    ff_ram[16111] = 8'h00;
    ff_ram[16112] = 8'h00;
    ff_ram[16113] = 8'h00;
    ff_ram[16114] = 8'h00;
    ff_ram[16115] = 8'h00;
    ff_ram[16116] = 8'h00;
    ff_ram[16117] = 8'h00;
    ff_ram[16118] = 8'h00;
    ff_ram[16119] = 8'h00;
    ff_ram[16120] = 8'h00;
    ff_ram[16121] = 8'h00;
    ff_ram[16122] = 8'h00;
    ff_ram[16123] = 8'h00;
    ff_ram[16124] = 8'h00;
    ff_ram[16125] = 8'h00;
    ff_ram[16126] = 8'h00;
    ff_ram[16127] = 8'h00;
    ff_ram[16128] = 8'h00;
    ff_ram[16129] = 8'h00;
    ff_ram[16130] = 8'h00;
    ff_ram[16131] = 8'h00;
    ff_ram[16132] = 8'h00;
    ff_ram[16133] = 8'h00;
    ff_ram[16134] = 8'h00;
    ff_ram[16135] = 8'h00;
    ff_ram[16136] = 8'h00;
    ff_ram[16137] = 8'h00;
    ff_ram[16138] = 8'h00;
    ff_ram[16139] = 8'h00;
    ff_ram[16140] = 8'h00;
    ff_ram[16141] = 8'h00;
    ff_ram[16142] = 8'h00;
    ff_ram[16143] = 8'h00;
    ff_ram[16144] = 8'h00;
    ff_ram[16145] = 8'h00;
    ff_ram[16146] = 8'h00;
    ff_ram[16147] = 8'h00;
    ff_ram[16148] = 8'h00;
    ff_ram[16149] = 8'h00;
    ff_ram[16150] = 8'h00;
    ff_ram[16151] = 8'h00;
    ff_ram[16152] = 8'h00;
    ff_ram[16153] = 8'h00;
    ff_ram[16154] = 8'h00;
    ff_ram[16155] = 8'h00;
    ff_ram[16156] = 8'h00;
    ff_ram[16157] = 8'h00;
    ff_ram[16158] = 8'h00;
    ff_ram[16159] = 8'h00;
    ff_ram[16160] = 8'h00;
    ff_ram[16161] = 8'h00;
    ff_ram[16162] = 8'h00;
    ff_ram[16163] = 8'h00;
    ff_ram[16164] = 8'h00;
    ff_ram[16165] = 8'h00;
    ff_ram[16166] = 8'h00;
    ff_ram[16167] = 8'h00;
    ff_ram[16168] = 8'h00;
    ff_ram[16169] = 8'h00;
    ff_ram[16170] = 8'h00;
    ff_ram[16171] = 8'h00;
    ff_ram[16172] = 8'h00;
    ff_ram[16173] = 8'h00;
    ff_ram[16174] = 8'h00;
    ff_ram[16175] = 8'h00;
    ff_ram[16176] = 8'h00;
    ff_ram[16177] = 8'h00;
    ff_ram[16178] = 8'h00;
    ff_ram[16179] = 8'h00;
    ff_ram[16180] = 8'h00;
    ff_ram[16181] = 8'h00;
    ff_ram[16182] = 8'h00;
    ff_ram[16183] = 8'h00;
    ff_ram[16184] = 8'h00;
    ff_ram[16185] = 8'h00;
    ff_ram[16186] = 8'h00;
    ff_ram[16187] = 8'h00;
    ff_ram[16188] = 8'h00;
    ff_ram[16189] = 8'h00;
    ff_ram[16190] = 8'h00;
    ff_ram[16191] = 8'h00;
    ff_ram[16192] = 8'h00;
    ff_ram[16193] = 8'h00;
    ff_ram[16194] = 8'h00;
    ff_ram[16195] = 8'h00;
    ff_ram[16196] = 8'h00;
    ff_ram[16197] = 8'h00;
    ff_ram[16198] = 8'h00;
    ff_ram[16199] = 8'h00;
    ff_ram[16200] = 8'h00;
    ff_ram[16201] = 8'h00;
    ff_ram[16202] = 8'h00;
    ff_ram[16203] = 8'h00;
    ff_ram[16204] = 8'h00;
    ff_ram[16205] = 8'h00;
    ff_ram[16206] = 8'h00;
    ff_ram[16207] = 8'h00;
    ff_ram[16208] = 8'h00;
    ff_ram[16209] = 8'h00;
    ff_ram[16210] = 8'h00;
    ff_ram[16211] = 8'h00;
    ff_ram[16212] = 8'h00;
    ff_ram[16213] = 8'h00;
    ff_ram[16214] = 8'h00;
    ff_ram[16215] = 8'h00;
    ff_ram[16216] = 8'h00;
    ff_ram[16217] = 8'h00;
    ff_ram[16218] = 8'h00;
    ff_ram[16219] = 8'h00;
    ff_ram[16220] = 8'h00;
    ff_ram[16221] = 8'h00;
    ff_ram[16222] = 8'h00;
    ff_ram[16223] = 8'h00;
    ff_ram[16224] = 8'h00;
    ff_ram[16225] = 8'h00;
    ff_ram[16226] = 8'h00;
    ff_ram[16227] = 8'h00;
    ff_ram[16228] = 8'h00;
    ff_ram[16229] = 8'h00;
    ff_ram[16230] = 8'h00;
    ff_ram[16231] = 8'h00;
    ff_ram[16232] = 8'h00;
    ff_ram[16233] = 8'h00;
    ff_ram[16234] = 8'h00;
    ff_ram[16235] = 8'h00;
    ff_ram[16236] = 8'h00;
    ff_ram[16237] = 8'h00;
    ff_ram[16238] = 8'h00;
    ff_ram[16239] = 8'h00;
    ff_ram[16240] = 8'h00;
    ff_ram[16241] = 8'h00;
    ff_ram[16242] = 8'h00;
    ff_ram[16243] = 8'h00;
    ff_ram[16244] = 8'h00;
    ff_ram[16245] = 8'h00;
    ff_ram[16246] = 8'h00;
    ff_ram[16247] = 8'h00;
    ff_ram[16248] = 8'h00;
    ff_ram[16249] = 8'h00;
    ff_ram[16250] = 8'h00;
    ff_ram[16251] = 8'h00;
    ff_ram[16252] = 8'h00;
    ff_ram[16253] = 8'h00;
    ff_ram[16254] = 8'h00;
    ff_ram[16255] = 8'h00;
    ff_ram[16256] = 8'h00;
    ff_ram[16257] = 8'h00;
    ff_ram[16258] = 8'h00;
    ff_ram[16259] = 8'h00;
    ff_ram[16260] = 8'h00;
    ff_ram[16261] = 8'h00;
    ff_ram[16262] = 8'h00;
    ff_ram[16263] = 8'h00;
    ff_ram[16264] = 8'h00;
    ff_ram[16265] = 8'h00;
    ff_ram[16266] = 8'h00;
    ff_ram[16267] = 8'h00;
    ff_ram[16268] = 8'h00;
    ff_ram[16269] = 8'h00;
    ff_ram[16270] = 8'h00;
    ff_ram[16271] = 8'h00;
    ff_ram[16272] = 8'h00;
    ff_ram[16273] = 8'h00;
    ff_ram[16274] = 8'h00;
    ff_ram[16275] = 8'h00;
    ff_ram[16276] = 8'h00;
    ff_ram[16277] = 8'h00;
    ff_ram[16278] = 8'h00;
    ff_ram[16279] = 8'h00;
    ff_ram[16280] = 8'h00;
    ff_ram[16281] = 8'h00;
    ff_ram[16282] = 8'h00;
    ff_ram[16283] = 8'h00;
    ff_ram[16284] = 8'h00;
    ff_ram[16285] = 8'h00;
    ff_ram[16286] = 8'h00;
    ff_ram[16287] = 8'h00;
    ff_ram[16288] = 8'h00;
    ff_ram[16289] = 8'h00;
    ff_ram[16290] = 8'h00;
    ff_ram[16291] = 8'h00;
    ff_ram[16292] = 8'h00;
    ff_ram[16293] = 8'h00;
    ff_ram[16294] = 8'h00;
    ff_ram[16295] = 8'h00;
    ff_ram[16296] = 8'h00;
    ff_ram[16297] = 8'h00;
    ff_ram[16298] = 8'h00;
    ff_ram[16299] = 8'h00;
    ff_ram[16300] = 8'h00;
    ff_ram[16301] = 8'h00;
    ff_ram[16302] = 8'h00;
    ff_ram[16303] = 8'h00;
    ff_ram[16304] = 8'h00;
    ff_ram[16305] = 8'h00;
    ff_ram[16306] = 8'h00;
    ff_ram[16307] = 8'h00;
    ff_ram[16308] = 8'h00;
    ff_ram[16309] = 8'h00;
    ff_ram[16310] = 8'h00;
    ff_ram[16311] = 8'h00;
    ff_ram[16312] = 8'h00;
    ff_ram[16313] = 8'h00;
    ff_ram[16314] = 8'h00;
    ff_ram[16315] = 8'h00;
    ff_ram[16316] = 8'h00;
    ff_ram[16317] = 8'h00;
    ff_ram[16318] = 8'h00;
    ff_ram[16319] = 8'h00;
    ff_ram[16320] = 8'h00;
    ff_ram[16321] = 8'h00;
    ff_ram[16322] = 8'h00;
    ff_ram[16323] = 8'h00;
    ff_ram[16324] = 8'h00;
    ff_ram[16325] = 8'h00;
    ff_ram[16326] = 8'h00;
    ff_ram[16327] = 8'h00;
    ff_ram[16328] = 8'h00;
    ff_ram[16329] = 8'h00;
    ff_ram[16330] = 8'h00;
    ff_ram[16331] = 8'h00;
    ff_ram[16332] = 8'h00;
    ff_ram[16333] = 8'h00;
    ff_ram[16334] = 8'h00;
    ff_ram[16335] = 8'h00;
    ff_ram[16336] = 8'h00;
    ff_ram[16337] = 8'h00;
    ff_ram[16338] = 8'h00;
    ff_ram[16339] = 8'h00;
    ff_ram[16340] = 8'h00;
    ff_ram[16341] = 8'h00;
    ff_ram[16342] = 8'h00;
    ff_ram[16343] = 8'h00;
    ff_ram[16344] = 8'h00;
    ff_ram[16345] = 8'h00;
    ff_ram[16346] = 8'h00;
    ff_ram[16347] = 8'h00;
    ff_ram[16348] = 8'h00;
    ff_ram[16349] = 8'h00;
    ff_ram[16350] = 8'h00;
    ff_ram[16351] = 8'h00;
    ff_ram[16352] = 8'h00;
    ff_ram[16353] = 8'h00;
    ff_ram[16354] = 8'h00;
    ff_ram[16355] = 8'h00;
    ff_ram[16356] = 8'h00;
    ff_ram[16357] = 8'h00;
    ff_ram[16358] = 8'h00;
    ff_ram[16359] = 8'h00;
    ff_ram[16360] = 8'h00;
    ff_ram[16361] = 8'h00;
    ff_ram[16362] = 8'h00;
    ff_ram[16363] = 8'h00;
    ff_ram[16364] = 8'h00;
    ff_ram[16365] = 8'h00;
    ff_ram[16366] = 8'h00;
    ff_ram[16367] = 8'h00;
    ff_ram[16368] = 8'h00;
    ff_ram[16369] = 8'h00;
    ff_ram[16370] = 8'h00;
    ff_ram[16371] = 8'h00;
    ff_ram[16372] = 8'h00;
    ff_ram[16373] = 8'h00;
    ff_ram[16374] = 8'h00;
    ff_ram[16375] = 8'h00;
    ff_ram[16376] = 8'h00;
    ff_ram[16377] = 8'h00;
    ff_ram[16378] = 8'h00;
    ff_ram[16379] = 8'h00;
    ff_ram[16380] = 8'h00;
    ff_ram[16381] = 8'h00;
    ff_ram[16382] = 8'h00;
    ff_ram[16383] = 8'h00;
end
