module Gowin_PLL(
	output			clkout,
	input			clkin
);
	assign clkout = clkin;
endmodule
