// romfont.bin���玩���������ꂽSystemVerilog�R�[�h
// ��������: 2025-08-11 21:06:54.461605

write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h54 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h12 );
write_io( vdp_io0, 8'h14 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h14 );
write_io( vdp_io0, 8'h34 );
write_io( vdp_io0, 8'h52 );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h54 );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h54 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h3C );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h86 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'hEE );
write_io( vdp_io0, 8'hA4 );
write_io( vdp_io0, 8'hEF );
write_io( vdp_io0, 8'hA2 );
write_io( vdp_io0, 8'hEA );
write_io( vdp_io0, 8'h06 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h3C );
write_io( vdp_io0, 8'h14 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h4C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h5C );
write_io( vdp_io0, 8'hEA );
write_io( vdp_io0, 8'h6C );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h0C );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h1E );
write_io( vdp_io0, 8'h12 );
write_io( vdp_io0, 8'h22 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h4E );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFF );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hFF );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h1F );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFF );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hFF );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h1F );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h1F );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h81 );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'h81 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h54 );
write_io( vdp_io0, 8'h54 );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hB8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hD8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hD8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hB0 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'hB0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hD0 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hB0 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hB0 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'hB0 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hB0 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h6C );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'hD6 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h4C );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h3C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'hB4 );
write_io( vdp_io0, 8'h64 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'hA4 );
write_io( vdp_io0, 8'h68 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h58 );
write_io( vdp_io0, 8'h64 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hB8 );
write_io( vdp_io0, 8'hD4 );
write_io( vdp_io0, 8'h94 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h1C );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h74 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'hAA );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h64 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h82 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h9C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'hFA );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'hA2 );
write_io( vdp_io0, 8'hA2 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'hF2 );
write_io( vdp_io0, 8'h4A );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h9E );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h3C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h3C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h28 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hC8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hD0 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'hE8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hA0 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'hA8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF0 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h58 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hC0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hE0 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h4E );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h8E );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'h02 );
write_io( vdp_io0, 8'h02 );
write_io( vdp_io0, 8'h02 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'hFE );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h1C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h2C );
write_io( vdp_io0, 8'hF2 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h9C );
write_io( vdp_io0, 8'h26 );
write_io( vdp_io0, 8'h1C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h9E );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'h90 );
write_io( vdp_io0, 8'h4E );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'hD2 );
write_io( vdp_io0, 8'hB6 );
write_io( vdp_io0, 8'hAA );
write_io( vdp_io0, 8'h4C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h4C );
write_io( vdp_io0, 8'hD2 );
write_io( vdp_io0, 8'h62 );
write_io( vdp_io0, 8'h4E );
write_io( vdp_io0, 8'hD2 );
write_io( vdp_io0, 8'h4E );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h54 );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'hA2 );
write_io( vdp_io0, 8'hA2 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h9E );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h8C );
write_io( vdp_io0, 8'h96 );
write_io( vdp_io0, 8'h4C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hE4 );
write_io( vdp_io0, 8'h26 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h14 );
write_io( vdp_io0, 8'h52 );
write_io( vdp_io0, 8'hB2 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h50 );
write_io( vdp_io0, 8'h88 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h02 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h1E );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h9E );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h8C );
write_io( vdp_io0, 8'h96 );
write_io( vdp_io0, 8'h4C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'hFC );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h98 );
write_io( vdp_io0, 8'h74 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h14 );
write_io( vdp_io0, 8'h7E );
write_io( vdp_io0, 8'hA4 );
write_io( vdp_io0, 8'hA4 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF4 );
write_io( vdp_io0, 8'h22 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'hA2 );
write_io( vdp_io0, 8'h62 );
write_io( vdp_io0, 8'h1C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h7C );
write_io( vdp_io0, 8'hAA );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'hA2 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'hF8 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h18 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h48 );
write_io( vdp_io0, 8'h5C );
write_io( vdp_io0, 8'h6A );
write_io( vdp_io0, 8'hE2 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h9C );
write_io( vdp_io0, 8'hB2 );
write_io( vdp_io0, 8'hD2 );
write_io( vdp_io0, 8'h92 );
write_io( vdp_io0, 8'h1C );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h1C );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h94 );
write_io( vdp_io0, 8'h70 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h80 );
write_io( vdp_io0, 8'hB8 );
write_io( vdp_io0, 8'hC4 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h08 );
write_io( vdp_io0, 8'h30 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'hB4 );
write_io( vdp_io0, 8'h4C );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h2C );
write_io( vdp_io0, 8'hF4 );
write_io( vdp_io0, 8'h24 );
write_io( vdp_io0, 8'h64 );
write_io( vdp_io0, 8'hA4 );
write_io( vdp_io0, 8'h26 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h78 );
write_io( vdp_io0, 8'h84 );
write_io( vdp_io0, 8'h04 );
write_io( vdp_io0, 8'h38 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'h40 );
write_io( vdp_io0, 8'hDC );
write_io( vdp_io0, 8'h62 );
write_io( vdp_io0, 8'h42 );
write_io( vdp_io0, 8'hC2 );
write_io( vdp_io0, 8'h44 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h10 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h20 );
write_io( vdp_io0, 8'h60 );
write_io( vdp_io0, 8'h52 );
write_io( vdp_io0, 8'h8C );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
write_io( vdp_io0, 8'h00 );
